`timescale 1 ns/100 ps
// Version: 2023.2 2023.2.0.8


module PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM(
       A_DIN,
       A_DOUT,
       B_DIN,
       B_DOUT,
       A_ADDR,
       B_ADDR,
       B_BLK_EN,
       A_REN,
       A_CLK,
       B_CLK,
       A_WEN,
       B_WEN,
       A_WBYTE_EN,
       B_WBYTE_EN
    );
input  [39:0] A_DIN;
output [39:0] A_DOUT;
input  [39:0] B_DIN;
output [39:0] B_DOUT;
input  [18:0] A_ADDR;
input  [18:0] B_ADDR;
input  B_BLK_EN;
input  A_REN;
input  A_CLK;
input  B_CLK;
input  A_WEN;
input  B_WEN;
input  [7:0] A_WBYTE_EN;
input  [7:0] B_WBYTE_EN;

    wire \WBYTEENA[0] , \WBYTEENA[2] , \WBYTEENA[4] , \WBYTEENA[6] , 
        \WBYTEENA[8] , \WBYTEENA[10] , \WBYTEENA[12] , \WBYTEENA[14] , 
        \WBYTEENB[0] , \WBYTEENB[2] , \WBYTEENB[4] , \WBYTEENB[6] , 
        \WBYTEENB[8] , \WBYTEENB[10] , \WBYTEENB[12] , \WBYTEENB[14] , 
        \B_DOUT_TEMPR0[0] , \B_DOUT_TEMPR1[0] , \B_DOUT_TEMPR2[0] , 
        \B_DOUT_TEMPR3[0] , \B_DOUT_TEMPR4[0] , \B_DOUT_TEMPR5[0] , 
        \B_DOUT_TEMPR6[0] , \B_DOUT_TEMPR7[0] , \B_DOUT_TEMPR8[0] , 
        \B_DOUT_TEMPR9[0] , \B_DOUT_TEMPR10[0] , \B_DOUT_TEMPR11[0] , 
        \B_DOUT_TEMPR12[0] , \B_DOUT_TEMPR13[0] , \B_DOUT_TEMPR14[0] , 
        \B_DOUT_TEMPR15[0] , \B_DOUT_TEMPR16[0] , \B_DOUT_TEMPR17[0] , 
        \B_DOUT_TEMPR18[0] , \B_DOUT_TEMPR19[0] , \B_DOUT_TEMPR20[0] , 
        \B_DOUT_TEMPR21[0] , \B_DOUT_TEMPR22[0] , \B_DOUT_TEMPR23[0] , 
        \B_DOUT_TEMPR24[0] , \B_DOUT_TEMPR25[0] , \B_DOUT_TEMPR26[0] , 
        \B_DOUT_TEMPR27[0] , \B_DOUT_TEMPR28[0] , \B_DOUT_TEMPR29[0] , 
        \B_DOUT_TEMPR30[0] , \B_DOUT_TEMPR31[0] , \B_DOUT_TEMPR32[0] , 
        \B_DOUT_TEMPR33[0] , \B_DOUT_TEMPR34[0] , \B_DOUT_TEMPR35[0] , 
        \B_DOUT_TEMPR36[0] , \B_DOUT_TEMPR37[0] , \B_DOUT_TEMPR38[0] , 
        \B_DOUT_TEMPR39[0] , \B_DOUT_TEMPR40[0] , \B_DOUT_TEMPR41[0] , 
        \B_DOUT_TEMPR42[0] , \B_DOUT_TEMPR43[0] , \B_DOUT_TEMPR44[0] , 
        \B_DOUT_TEMPR45[0] , \B_DOUT_TEMPR46[0] , \B_DOUT_TEMPR47[0] , 
        \B_DOUT_TEMPR48[0] , \B_DOUT_TEMPR49[0] , \B_DOUT_TEMPR50[0] , 
        \B_DOUT_TEMPR51[0] , \B_DOUT_TEMPR52[0] , \B_DOUT_TEMPR53[0] , 
        \B_DOUT_TEMPR54[0] , \B_DOUT_TEMPR55[0] , \B_DOUT_TEMPR56[0] , 
        \B_DOUT_TEMPR57[0] , \B_DOUT_TEMPR58[0] , \B_DOUT_TEMPR59[0] , 
        \B_DOUT_TEMPR60[0] , \B_DOUT_TEMPR61[0] , \B_DOUT_TEMPR62[0] , 
        \B_DOUT_TEMPR63[0] , \B_DOUT_TEMPR64[0] , \B_DOUT_TEMPR65[0] , 
        \B_DOUT_TEMPR66[0] , \B_DOUT_TEMPR67[0] , \B_DOUT_TEMPR68[0] , 
        \B_DOUT_TEMPR69[0] , \B_DOUT_TEMPR70[0] , \B_DOUT_TEMPR71[0] , 
        \B_DOUT_TEMPR72[0] , \B_DOUT_TEMPR73[0] , \B_DOUT_TEMPR74[0] , 
        \B_DOUT_TEMPR75[0] , \B_DOUT_TEMPR76[0] , \B_DOUT_TEMPR77[0] , 
        \B_DOUT_TEMPR78[0] , \B_DOUT_TEMPR79[0] , \B_DOUT_TEMPR80[0] , 
        \B_DOUT_TEMPR81[0] , \B_DOUT_TEMPR82[0] , \B_DOUT_TEMPR83[0] , 
        \B_DOUT_TEMPR84[0] , \B_DOUT_TEMPR85[0] , \B_DOUT_TEMPR86[0] , 
        \B_DOUT_TEMPR87[0] , \B_DOUT_TEMPR88[0] , \B_DOUT_TEMPR89[0] , 
        \B_DOUT_TEMPR90[0] , \B_DOUT_TEMPR91[0] , \B_DOUT_TEMPR92[0] , 
        \B_DOUT_TEMPR93[0] , \B_DOUT_TEMPR94[0] , \B_DOUT_TEMPR95[0] , 
        \B_DOUT_TEMPR96[0] , \B_DOUT_TEMPR97[0] , \B_DOUT_TEMPR98[0] , 
        \B_DOUT_TEMPR99[0] , \B_DOUT_TEMPR100[0] , 
        \B_DOUT_TEMPR101[0] , \B_DOUT_TEMPR102[0] , 
        \B_DOUT_TEMPR103[0] , \B_DOUT_TEMPR104[0] , 
        \B_DOUT_TEMPR105[0] , \B_DOUT_TEMPR106[0] , 
        \B_DOUT_TEMPR107[0] , \B_DOUT_TEMPR108[0] , 
        \B_DOUT_TEMPR109[0] , \B_DOUT_TEMPR110[0] , 
        \B_DOUT_TEMPR111[0] , \B_DOUT_TEMPR112[0] , 
        \B_DOUT_TEMPR113[0] , \B_DOUT_TEMPR114[0] , 
        \B_DOUT_TEMPR115[0] , \B_DOUT_TEMPR116[0] , 
        \B_DOUT_TEMPR117[0] , \B_DOUT_TEMPR118[0] , \B_DOUT_TEMPR0[1] , 
        \B_DOUT_TEMPR1[1] , \B_DOUT_TEMPR2[1] , \B_DOUT_TEMPR3[1] , 
        \B_DOUT_TEMPR4[1] , \B_DOUT_TEMPR5[1] , \B_DOUT_TEMPR6[1] , 
        \B_DOUT_TEMPR7[1] , \B_DOUT_TEMPR8[1] , \B_DOUT_TEMPR9[1] , 
        \B_DOUT_TEMPR10[1] , \B_DOUT_TEMPR11[1] , \B_DOUT_TEMPR12[1] , 
        \B_DOUT_TEMPR13[1] , \B_DOUT_TEMPR14[1] , \B_DOUT_TEMPR15[1] , 
        \B_DOUT_TEMPR16[1] , \B_DOUT_TEMPR17[1] , \B_DOUT_TEMPR18[1] , 
        \B_DOUT_TEMPR19[1] , \B_DOUT_TEMPR20[1] , \B_DOUT_TEMPR21[1] , 
        \B_DOUT_TEMPR22[1] , \B_DOUT_TEMPR23[1] , \B_DOUT_TEMPR24[1] , 
        \B_DOUT_TEMPR25[1] , \B_DOUT_TEMPR26[1] , \B_DOUT_TEMPR27[1] , 
        \B_DOUT_TEMPR28[1] , \B_DOUT_TEMPR29[1] , \B_DOUT_TEMPR30[1] , 
        \B_DOUT_TEMPR31[1] , \B_DOUT_TEMPR32[1] , \B_DOUT_TEMPR33[1] , 
        \B_DOUT_TEMPR34[1] , \B_DOUT_TEMPR35[1] , \B_DOUT_TEMPR36[1] , 
        \B_DOUT_TEMPR37[1] , \B_DOUT_TEMPR38[1] , \B_DOUT_TEMPR39[1] , 
        \B_DOUT_TEMPR40[1] , \B_DOUT_TEMPR41[1] , \B_DOUT_TEMPR42[1] , 
        \B_DOUT_TEMPR43[1] , \B_DOUT_TEMPR44[1] , \B_DOUT_TEMPR45[1] , 
        \B_DOUT_TEMPR46[1] , \B_DOUT_TEMPR47[1] , \B_DOUT_TEMPR48[1] , 
        \B_DOUT_TEMPR49[1] , \B_DOUT_TEMPR50[1] , \B_DOUT_TEMPR51[1] , 
        \B_DOUT_TEMPR52[1] , \B_DOUT_TEMPR53[1] , \B_DOUT_TEMPR54[1] , 
        \B_DOUT_TEMPR55[1] , \B_DOUT_TEMPR56[1] , \B_DOUT_TEMPR57[1] , 
        \B_DOUT_TEMPR58[1] , \B_DOUT_TEMPR59[1] , \B_DOUT_TEMPR60[1] , 
        \B_DOUT_TEMPR61[1] , \B_DOUT_TEMPR62[1] , \B_DOUT_TEMPR63[1] , 
        \B_DOUT_TEMPR64[1] , \B_DOUT_TEMPR65[1] , \B_DOUT_TEMPR66[1] , 
        \B_DOUT_TEMPR67[1] , \B_DOUT_TEMPR68[1] , \B_DOUT_TEMPR69[1] , 
        \B_DOUT_TEMPR70[1] , \B_DOUT_TEMPR71[1] , \B_DOUT_TEMPR72[1] , 
        \B_DOUT_TEMPR73[1] , \B_DOUT_TEMPR74[1] , \B_DOUT_TEMPR75[1] , 
        \B_DOUT_TEMPR76[1] , \B_DOUT_TEMPR77[1] , \B_DOUT_TEMPR78[1] , 
        \B_DOUT_TEMPR79[1] , \B_DOUT_TEMPR80[1] , \B_DOUT_TEMPR81[1] , 
        \B_DOUT_TEMPR82[1] , \B_DOUT_TEMPR83[1] , \B_DOUT_TEMPR84[1] , 
        \B_DOUT_TEMPR85[1] , \B_DOUT_TEMPR86[1] , \B_DOUT_TEMPR87[1] , 
        \B_DOUT_TEMPR88[1] , \B_DOUT_TEMPR89[1] , \B_DOUT_TEMPR90[1] , 
        \B_DOUT_TEMPR91[1] , \B_DOUT_TEMPR92[1] , \B_DOUT_TEMPR93[1] , 
        \B_DOUT_TEMPR94[1] , \B_DOUT_TEMPR95[1] , \B_DOUT_TEMPR96[1] , 
        \B_DOUT_TEMPR97[1] , \B_DOUT_TEMPR98[1] , \B_DOUT_TEMPR99[1] , 
        \B_DOUT_TEMPR100[1] , \B_DOUT_TEMPR101[1] , 
        \B_DOUT_TEMPR102[1] , \B_DOUT_TEMPR103[1] , 
        \B_DOUT_TEMPR104[1] , \B_DOUT_TEMPR105[1] , 
        \B_DOUT_TEMPR106[1] , \B_DOUT_TEMPR107[1] , 
        \B_DOUT_TEMPR108[1] , \B_DOUT_TEMPR109[1] , 
        \B_DOUT_TEMPR110[1] , \B_DOUT_TEMPR111[1] , 
        \B_DOUT_TEMPR112[1] , \B_DOUT_TEMPR113[1] , 
        \B_DOUT_TEMPR114[1] , \B_DOUT_TEMPR115[1] , 
        \B_DOUT_TEMPR116[1] , \B_DOUT_TEMPR117[1] , 
        \B_DOUT_TEMPR118[1] , \B_DOUT_TEMPR0[2] , \B_DOUT_TEMPR1[2] , 
        \B_DOUT_TEMPR2[2] , \B_DOUT_TEMPR3[2] , \B_DOUT_TEMPR4[2] , 
        \B_DOUT_TEMPR5[2] , \B_DOUT_TEMPR6[2] , \B_DOUT_TEMPR7[2] , 
        \B_DOUT_TEMPR8[2] , \B_DOUT_TEMPR9[2] , \B_DOUT_TEMPR10[2] , 
        \B_DOUT_TEMPR11[2] , \B_DOUT_TEMPR12[2] , \B_DOUT_TEMPR13[2] , 
        \B_DOUT_TEMPR14[2] , \B_DOUT_TEMPR15[2] , \B_DOUT_TEMPR16[2] , 
        \B_DOUT_TEMPR17[2] , \B_DOUT_TEMPR18[2] , \B_DOUT_TEMPR19[2] , 
        \B_DOUT_TEMPR20[2] , \B_DOUT_TEMPR21[2] , \B_DOUT_TEMPR22[2] , 
        \B_DOUT_TEMPR23[2] , \B_DOUT_TEMPR24[2] , \B_DOUT_TEMPR25[2] , 
        \B_DOUT_TEMPR26[2] , \B_DOUT_TEMPR27[2] , \B_DOUT_TEMPR28[2] , 
        \B_DOUT_TEMPR29[2] , \B_DOUT_TEMPR30[2] , \B_DOUT_TEMPR31[2] , 
        \B_DOUT_TEMPR32[2] , \B_DOUT_TEMPR33[2] , \B_DOUT_TEMPR34[2] , 
        \B_DOUT_TEMPR35[2] , \B_DOUT_TEMPR36[2] , \B_DOUT_TEMPR37[2] , 
        \B_DOUT_TEMPR38[2] , \B_DOUT_TEMPR39[2] , \B_DOUT_TEMPR40[2] , 
        \B_DOUT_TEMPR41[2] , \B_DOUT_TEMPR42[2] , \B_DOUT_TEMPR43[2] , 
        \B_DOUT_TEMPR44[2] , \B_DOUT_TEMPR45[2] , \B_DOUT_TEMPR46[2] , 
        \B_DOUT_TEMPR47[2] , \B_DOUT_TEMPR48[2] , \B_DOUT_TEMPR49[2] , 
        \B_DOUT_TEMPR50[2] , \B_DOUT_TEMPR51[2] , \B_DOUT_TEMPR52[2] , 
        \B_DOUT_TEMPR53[2] , \B_DOUT_TEMPR54[2] , \B_DOUT_TEMPR55[2] , 
        \B_DOUT_TEMPR56[2] , \B_DOUT_TEMPR57[2] , \B_DOUT_TEMPR58[2] , 
        \B_DOUT_TEMPR59[2] , \B_DOUT_TEMPR60[2] , \B_DOUT_TEMPR61[2] , 
        \B_DOUT_TEMPR62[2] , \B_DOUT_TEMPR63[2] , \B_DOUT_TEMPR64[2] , 
        \B_DOUT_TEMPR65[2] , \B_DOUT_TEMPR66[2] , \B_DOUT_TEMPR67[2] , 
        \B_DOUT_TEMPR68[2] , \B_DOUT_TEMPR69[2] , \B_DOUT_TEMPR70[2] , 
        \B_DOUT_TEMPR71[2] , \B_DOUT_TEMPR72[2] , \B_DOUT_TEMPR73[2] , 
        \B_DOUT_TEMPR74[2] , \B_DOUT_TEMPR75[2] , \B_DOUT_TEMPR76[2] , 
        \B_DOUT_TEMPR77[2] , \B_DOUT_TEMPR78[2] , \B_DOUT_TEMPR79[2] , 
        \B_DOUT_TEMPR80[2] , \B_DOUT_TEMPR81[2] , \B_DOUT_TEMPR82[2] , 
        \B_DOUT_TEMPR83[2] , \B_DOUT_TEMPR84[2] , \B_DOUT_TEMPR85[2] , 
        \B_DOUT_TEMPR86[2] , \B_DOUT_TEMPR87[2] , \B_DOUT_TEMPR88[2] , 
        \B_DOUT_TEMPR89[2] , \B_DOUT_TEMPR90[2] , \B_DOUT_TEMPR91[2] , 
        \B_DOUT_TEMPR92[2] , \B_DOUT_TEMPR93[2] , \B_DOUT_TEMPR94[2] , 
        \B_DOUT_TEMPR95[2] , \B_DOUT_TEMPR96[2] , \B_DOUT_TEMPR97[2] , 
        \B_DOUT_TEMPR98[2] , \B_DOUT_TEMPR99[2] , \B_DOUT_TEMPR100[2] , 
        \B_DOUT_TEMPR101[2] , \B_DOUT_TEMPR102[2] , 
        \B_DOUT_TEMPR103[2] , \B_DOUT_TEMPR104[2] , 
        \B_DOUT_TEMPR105[2] , \B_DOUT_TEMPR106[2] , 
        \B_DOUT_TEMPR107[2] , \B_DOUT_TEMPR108[2] , 
        \B_DOUT_TEMPR109[2] , \B_DOUT_TEMPR110[2] , 
        \B_DOUT_TEMPR111[2] , \B_DOUT_TEMPR112[2] , 
        \B_DOUT_TEMPR113[2] , \B_DOUT_TEMPR114[2] , 
        \B_DOUT_TEMPR115[2] , \B_DOUT_TEMPR116[2] , 
        \B_DOUT_TEMPR117[2] , \B_DOUT_TEMPR118[2] , \B_DOUT_TEMPR0[3] , 
        \B_DOUT_TEMPR1[3] , \B_DOUT_TEMPR2[3] , \B_DOUT_TEMPR3[3] , 
        \B_DOUT_TEMPR4[3] , \B_DOUT_TEMPR5[3] , \B_DOUT_TEMPR6[3] , 
        \B_DOUT_TEMPR7[3] , \B_DOUT_TEMPR8[3] , \B_DOUT_TEMPR9[3] , 
        \B_DOUT_TEMPR10[3] , \B_DOUT_TEMPR11[3] , \B_DOUT_TEMPR12[3] , 
        \B_DOUT_TEMPR13[3] , \B_DOUT_TEMPR14[3] , \B_DOUT_TEMPR15[3] , 
        \B_DOUT_TEMPR16[3] , \B_DOUT_TEMPR17[3] , \B_DOUT_TEMPR18[3] , 
        \B_DOUT_TEMPR19[3] , \B_DOUT_TEMPR20[3] , \B_DOUT_TEMPR21[3] , 
        \B_DOUT_TEMPR22[3] , \B_DOUT_TEMPR23[3] , \B_DOUT_TEMPR24[3] , 
        \B_DOUT_TEMPR25[3] , \B_DOUT_TEMPR26[3] , \B_DOUT_TEMPR27[3] , 
        \B_DOUT_TEMPR28[3] , \B_DOUT_TEMPR29[3] , \B_DOUT_TEMPR30[3] , 
        \B_DOUT_TEMPR31[3] , \B_DOUT_TEMPR32[3] , \B_DOUT_TEMPR33[3] , 
        \B_DOUT_TEMPR34[3] , \B_DOUT_TEMPR35[3] , \B_DOUT_TEMPR36[3] , 
        \B_DOUT_TEMPR37[3] , \B_DOUT_TEMPR38[3] , \B_DOUT_TEMPR39[3] , 
        \B_DOUT_TEMPR40[3] , \B_DOUT_TEMPR41[3] , \B_DOUT_TEMPR42[3] , 
        \B_DOUT_TEMPR43[3] , \B_DOUT_TEMPR44[3] , \B_DOUT_TEMPR45[3] , 
        \B_DOUT_TEMPR46[3] , \B_DOUT_TEMPR47[3] , \B_DOUT_TEMPR48[3] , 
        \B_DOUT_TEMPR49[3] , \B_DOUT_TEMPR50[3] , \B_DOUT_TEMPR51[3] , 
        \B_DOUT_TEMPR52[3] , \B_DOUT_TEMPR53[3] , \B_DOUT_TEMPR54[3] , 
        \B_DOUT_TEMPR55[3] , \B_DOUT_TEMPR56[3] , \B_DOUT_TEMPR57[3] , 
        \B_DOUT_TEMPR58[3] , \B_DOUT_TEMPR59[3] , \B_DOUT_TEMPR60[3] , 
        \B_DOUT_TEMPR61[3] , \B_DOUT_TEMPR62[3] , \B_DOUT_TEMPR63[3] , 
        \B_DOUT_TEMPR64[3] , \B_DOUT_TEMPR65[3] , \B_DOUT_TEMPR66[3] , 
        \B_DOUT_TEMPR67[3] , \B_DOUT_TEMPR68[3] , \B_DOUT_TEMPR69[3] , 
        \B_DOUT_TEMPR70[3] , \B_DOUT_TEMPR71[3] , \B_DOUT_TEMPR72[3] , 
        \B_DOUT_TEMPR73[3] , \B_DOUT_TEMPR74[3] , \B_DOUT_TEMPR75[3] , 
        \B_DOUT_TEMPR76[3] , \B_DOUT_TEMPR77[3] , \B_DOUT_TEMPR78[3] , 
        \B_DOUT_TEMPR79[3] , \B_DOUT_TEMPR80[3] , \B_DOUT_TEMPR81[3] , 
        \B_DOUT_TEMPR82[3] , \B_DOUT_TEMPR83[3] , \B_DOUT_TEMPR84[3] , 
        \B_DOUT_TEMPR85[3] , \B_DOUT_TEMPR86[3] , \B_DOUT_TEMPR87[3] , 
        \B_DOUT_TEMPR88[3] , \B_DOUT_TEMPR89[3] , \B_DOUT_TEMPR90[3] , 
        \B_DOUT_TEMPR91[3] , \B_DOUT_TEMPR92[3] , \B_DOUT_TEMPR93[3] , 
        \B_DOUT_TEMPR94[3] , \B_DOUT_TEMPR95[3] , \B_DOUT_TEMPR96[3] , 
        \B_DOUT_TEMPR97[3] , \B_DOUT_TEMPR98[3] , \B_DOUT_TEMPR99[3] , 
        \B_DOUT_TEMPR100[3] , \B_DOUT_TEMPR101[3] , 
        \B_DOUT_TEMPR102[3] , \B_DOUT_TEMPR103[3] , 
        \B_DOUT_TEMPR104[3] , \B_DOUT_TEMPR105[3] , 
        \B_DOUT_TEMPR106[3] , \B_DOUT_TEMPR107[3] , 
        \B_DOUT_TEMPR108[3] , \B_DOUT_TEMPR109[3] , 
        \B_DOUT_TEMPR110[3] , \B_DOUT_TEMPR111[3] , 
        \B_DOUT_TEMPR112[3] , \B_DOUT_TEMPR113[3] , 
        \B_DOUT_TEMPR114[3] , \B_DOUT_TEMPR115[3] , 
        \B_DOUT_TEMPR116[3] , \B_DOUT_TEMPR117[3] , 
        \B_DOUT_TEMPR118[3] , \B_DOUT_TEMPR0[4] , \B_DOUT_TEMPR1[4] , 
        \B_DOUT_TEMPR2[4] , \B_DOUT_TEMPR3[4] , \B_DOUT_TEMPR4[4] , 
        \B_DOUT_TEMPR5[4] , \B_DOUT_TEMPR6[4] , \B_DOUT_TEMPR7[4] , 
        \B_DOUT_TEMPR8[4] , \B_DOUT_TEMPR9[4] , \B_DOUT_TEMPR10[4] , 
        \B_DOUT_TEMPR11[4] , \B_DOUT_TEMPR12[4] , \B_DOUT_TEMPR13[4] , 
        \B_DOUT_TEMPR14[4] , \B_DOUT_TEMPR15[4] , \B_DOUT_TEMPR16[4] , 
        \B_DOUT_TEMPR17[4] , \B_DOUT_TEMPR18[4] , \B_DOUT_TEMPR19[4] , 
        \B_DOUT_TEMPR20[4] , \B_DOUT_TEMPR21[4] , \B_DOUT_TEMPR22[4] , 
        \B_DOUT_TEMPR23[4] , \B_DOUT_TEMPR24[4] , \B_DOUT_TEMPR25[4] , 
        \B_DOUT_TEMPR26[4] , \B_DOUT_TEMPR27[4] , \B_DOUT_TEMPR28[4] , 
        \B_DOUT_TEMPR29[4] , \B_DOUT_TEMPR30[4] , \B_DOUT_TEMPR31[4] , 
        \B_DOUT_TEMPR32[4] , \B_DOUT_TEMPR33[4] , \B_DOUT_TEMPR34[4] , 
        \B_DOUT_TEMPR35[4] , \B_DOUT_TEMPR36[4] , \B_DOUT_TEMPR37[4] , 
        \B_DOUT_TEMPR38[4] , \B_DOUT_TEMPR39[4] , \B_DOUT_TEMPR40[4] , 
        \B_DOUT_TEMPR41[4] , \B_DOUT_TEMPR42[4] , \B_DOUT_TEMPR43[4] , 
        \B_DOUT_TEMPR44[4] , \B_DOUT_TEMPR45[4] , \B_DOUT_TEMPR46[4] , 
        \B_DOUT_TEMPR47[4] , \B_DOUT_TEMPR48[4] , \B_DOUT_TEMPR49[4] , 
        \B_DOUT_TEMPR50[4] , \B_DOUT_TEMPR51[4] , \B_DOUT_TEMPR52[4] , 
        \B_DOUT_TEMPR53[4] , \B_DOUT_TEMPR54[4] , \B_DOUT_TEMPR55[4] , 
        \B_DOUT_TEMPR56[4] , \B_DOUT_TEMPR57[4] , \B_DOUT_TEMPR58[4] , 
        \B_DOUT_TEMPR59[4] , \B_DOUT_TEMPR60[4] , \B_DOUT_TEMPR61[4] , 
        \B_DOUT_TEMPR62[4] , \B_DOUT_TEMPR63[4] , \B_DOUT_TEMPR64[4] , 
        \B_DOUT_TEMPR65[4] , \B_DOUT_TEMPR66[4] , \B_DOUT_TEMPR67[4] , 
        \B_DOUT_TEMPR68[4] , \B_DOUT_TEMPR69[4] , \B_DOUT_TEMPR70[4] , 
        \B_DOUT_TEMPR71[4] , \B_DOUT_TEMPR72[4] , \B_DOUT_TEMPR73[4] , 
        \B_DOUT_TEMPR74[4] , \B_DOUT_TEMPR75[4] , \B_DOUT_TEMPR76[4] , 
        \B_DOUT_TEMPR77[4] , \B_DOUT_TEMPR78[4] , \B_DOUT_TEMPR79[4] , 
        \B_DOUT_TEMPR80[4] , \B_DOUT_TEMPR81[4] , \B_DOUT_TEMPR82[4] , 
        \B_DOUT_TEMPR83[4] , \B_DOUT_TEMPR84[4] , \B_DOUT_TEMPR85[4] , 
        \B_DOUT_TEMPR86[4] , \B_DOUT_TEMPR87[4] , \B_DOUT_TEMPR88[4] , 
        \B_DOUT_TEMPR89[4] , \B_DOUT_TEMPR90[4] , \B_DOUT_TEMPR91[4] , 
        \B_DOUT_TEMPR92[4] , \B_DOUT_TEMPR93[4] , \B_DOUT_TEMPR94[4] , 
        \B_DOUT_TEMPR95[4] , \B_DOUT_TEMPR96[4] , \B_DOUT_TEMPR97[4] , 
        \B_DOUT_TEMPR98[4] , \B_DOUT_TEMPR99[4] , \B_DOUT_TEMPR100[4] , 
        \B_DOUT_TEMPR101[4] , \B_DOUT_TEMPR102[4] , 
        \B_DOUT_TEMPR103[4] , \B_DOUT_TEMPR104[4] , 
        \B_DOUT_TEMPR105[4] , \B_DOUT_TEMPR106[4] , 
        \B_DOUT_TEMPR107[4] , \B_DOUT_TEMPR108[4] , 
        \B_DOUT_TEMPR109[4] , \B_DOUT_TEMPR110[4] , 
        \B_DOUT_TEMPR111[4] , \B_DOUT_TEMPR112[4] , 
        \B_DOUT_TEMPR113[4] , \B_DOUT_TEMPR114[4] , 
        \B_DOUT_TEMPR115[4] , \B_DOUT_TEMPR116[4] , 
        \B_DOUT_TEMPR117[4] , \B_DOUT_TEMPR118[4] , \B_DOUT_TEMPR0[5] , 
        \B_DOUT_TEMPR1[5] , \B_DOUT_TEMPR2[5] , \B_DOUT_TEMPR3[5] , 
        \B_DOUT_TEMPR4[5] , \B_DOUT_TEMPR5[5] , \B_DOUT_TEMPR6[5] , 
        \B_DOUT_TEMPR7[5] , \B_DOUT_TEMPR8[5] , \B_DOUT_TEMPR9[5] , 
        \B_DOUT_TEMPR10[5] , \B_DOUT_TEMPR11[5] , \B_DOUT_TEMPR12[5] , 
        \B_DOUT_TEMPR13[5] , \B_DOUT_TEMPR14[5] , \B_DOUT_TEMPR15[5] , 
        \B_DOUT_TEMPR16[5] , \B_DOUT_TEMPR17[5] , \B_DOUT_TEMPR18[5] , 
        \B_DOUT_TEMPR19[5] , \B_DOUT_TEMPR20[5] , \B_DOUT_TEMPR21[5] , 
        \B_DOUT_TEMPR22[5] , \B_DOUT_TEMPR23[5] , \B_DOUT_TEMPR24[5] , 
        \B_DOUT_TEMPR25[5] , \B_DOUT_TEMPR26[5] , \B_DOUT_TEMPR27[5] , 
        \B_DOUT_TEMPR28[5] , \B_DOUT_TEMPR29[5] , \B_DOUT_TEMPR30[5] , 
        \B_DOUT_TEMPR31[5] , \B_DOUT_TEMPR32[5] , \B_DOUT_TEMPR33[5] , 
        \B_DOUT_TEMPR34[5] , \B_DOUT_TEMPR35[5] , \B_DOUT_TEMPR36[5] , 
        \B_DOUT_TEMPR37[5] , \B_DOUT_TEMPR38[5] , \B_DOUT_TEMPR39[5] , 
        \B_DOUT_TEMPR40[5] , \B_DOUT_TEMPR41[5] , \B_DOUT_TEMPR42[5] , 
        \B_DOUT_TEMPR43[5] , \B_DOUT_TEMPR44[5] , \B_DOUT_TEMPR45[5] , 
        \B_DOUT_TEMPR46[5] , \B_DOUT_TEMPR47[5] , \B_DOUT_TEMPR48[5] , 
        \B_DOUT_TEMPR49[5] , \B_DOUT_TEMPR50[5] , \B_DOUT_TEMPR51[5] , 
        \B_DOUT_TEMPR52[5] , \B_DOUT_TEMPR53[5] , \B_DOUT_TEMPR54[5] , 
        \B_DOUT_TEMPR55[5] , \B_DOUT_TEMPR56[5] , \B_DOUT_TEMPR57[5] , 
        \B_DOUT_TEMPR58[5] , \B_DOUT_TEMPR59[5] , \B_DOUT_TEMPR60[5] , 
        \B_DOUT_TEMPR61[5] , \B_DOUT_TEMPR62[5] , \B_DOUT_TEMPR63[5] , 
        \B_DOUT_TEMPR64[5] , \B_DOUT_TEMPR65[5] , \B_DOUT_TEMPR66[5] , 
        \B_DOUT_TEMPR67[5] , \B_DOUT_TEMPR68[5] , \B_DOUT_TEMPR69[5] , 
        \B_DOUT_TEMPR70[5] , \B_DOUT_TEMPR71[5] , \B_DOUT_TEMPR72[5] , 
        \B_DOUT_TEMPR73[5] , \B_DOUT_TEMPR74[5] , \B_DOUT_TEMPR75[5] , 
        \B_DOUT_TEMPR76[5] , \B_DOUT_TEMPR77[5] , \B_DOUT_TEMPR78[5] , 
        \B_DOUT_TEMPR79[5] , \B_DOUT_TEMPR80[5] , \B_DOUT_TEMPR81[5] , 
        \B_DOUT_TEMPR82[5] , \B_DOUT_TEMPR83[5] , \B_DOUT_TEMPR84[5] , 
        \B_DOUT_TEMPR85[5] , \B_DOUT_TEMPR86[5] , \B_DOUT_TEMPR87[5] , 
        \B_DOUT_TEMPR88[5] , \B_DOUT_TEMPR89[5] , \B_DOUT_TEMPR90[5] , 
        \B_DOUT_TEMPR91[5] , \B_DOUT_TEMPR92[5] , \B_DOUT_TEMPR93[5] , 
        \B_DOUT_TEMPR94[5] , \B_DOUT_TEMPR95[5] , \B_DOUT_TEMPR96[5] , 
        \B_DOUT_TEMPR97[5] , \B_DOUT_TEMPR98[5] , \B_DOUT_TEMPR99[5] , 
        \B_DOUT_TEMPR100[5] , \B_DOUT_TEMPR101[5] , 
        \B_DOUT_TEMPR102[5] , \B_DOUT_TEMPR103[5] , 
        \B_DOUT_TEMPR104[5] , \B_DOUT_TEMPR105[5] , 
        \B_DOUT_TEMPR106[5] , \B_DOUT_TEMPR107[5] , 
        \B_DOUT_TEMPR108[5] , \B_DOUT_TEMPR109[5] , 
        \B_DOUT_TEMPR110[5] , \B_DOUT_TEMPR111[5] , 
        \B_DOUT_TEMPR112[5] , \B_DOUT_TEMPR113[5] , 
        \B_DOUT_TEMPR114[5] , \B_DOUT_TEMPR115[5] , 
        \B_DOUT_TEMPR116[5] , \B_DOUT_TEMPR117[5] , 
        \B_DOUT_TEMPR118[5] , \B_DOUT_TEMPR0[6] , \B_DOUT_TEMPR1[6] , 
        \B_DOUT_TEMPR2[6] , \B_DOUT_TEMPR3[6] , \B_DOUT_TEMPR4[6] , 
        \B_DOUT_TEMPR5[6] , \B_DOUT_TEMPR6[6] , \B_DOUT_TEMPR7[6] , 
        \B_DOUT_TEMPR8[6] , \B_DOUT_TEMPR9[6] , \B_DOUT_TEMPR10[6] , 
        \B_DOUT_TEMPR11[6] , \B_DOUT_TEMPR12[6] , \B_DOUT_TEMPR13[6] , 
        \B_DOUT_TEMPR14[6] , \B_DOUT_TEMPR15[6] , \B_DOUT_TEMPR16[6] , 
        \B_DOUT_TEMPR17[6] , \B_DOUT_TEMPR18[6] , \B_DOUT_TEMPR19[6] , 
        \B_DOUT_TEMPR20[6] , \B_DOUT_TEMPR21[6] , \B_DOUT_TEMPR22[6] , 
        \B_DOUT_TEMPR23[6] , \B_DOUT_TEMPR24[6] , \B_DOUT_TEMPR25[6] , 
        \B_DOUT_TEMPR26[6] , \B_DOUT_TEMPR27[6] , \B_DOUT_TEMPR28[6] , 
        \B_DOUT_TEMPR29[6] , \B_DOUT_TEMPR30[6] , \B_DOUT_TEMPR31[6] , 
        \B_DOUT_TEMPR32[6] , \B_DOUT_TEMPR33[6] , \B_DOUT_TEMPR34[6] , 
        \B_DOUT_TEMPR35[6] , \B_DOUT_TEMPR36[6] , \B_DOUT_TEMPR37[6] , 
        \B_DOUT_TEMPR38[6] , \B_DOUT_TEMPR39[6] , \B_DOUT_TEMPR40[6] , 
        \B_DOUT_TEMPR41[6] , \B_DOUT_TEMPR42[6] , \B_DOUT_TEMPR43[6] , 
        \B_DOUT_TEMPR44[6] , \B_DOUT_TEMPR45[6] , \B_DOUT_TEMPR46[6] , 
        \B_DOUT_TEMPR47[6] , \B_DOUT_TEMPR48[6] , \B_DOUT_TEMPR49[6] , 
        \B_DOUT_TEMPR50[6] , \B_DOUT_TEMPR51[6] , \B_DOUT_TEMPR52[6] , 
        \B_DOUT_TEMPR53[6] , \B_DOUT_TEMPR54[6] , \B_DOUT_TEMPR55[6] , 
        \B_DOUT_TEMPR56[6] , \B_DOUT_TEMPR57[6] , \B_DOUT_TEMPR58[6] , 
        \B_DOUT_TEMPR59[6] , \B_DOUT_TEMPR60[6] , \B_DOUT_TEMPR61[6] , 
        \B_DOUT_TEMPR62[6] , \B_DOUT_TEMPR63[6] , \B_DOUT_TEMPR64[6] , 
        \B_DOUT_TEMPR65[6] , \B_DOUT_TEMPR66[6] , \B_DOUT_TEMPR67[6] , 
        \B_DOUT_TEMPR68[6] , \B_DOUT_TEMPR69[6] , \B_DOUT_TEMPR70[6] , 
        \B_DOUT_TEMPR71[6] , \B_DOUT_TEMPR72[6] , \B_DOUT_TEMPR73[6] , 
        \B_DOUT_TEMPR74[6] , \B_DOUT_TEMPR75[6] , \B_DOUT_TEMPR76[6] , 
        \B_DOUT_TEMPR77[6] , \B_DOUT_TEMPR78[6] , \B_DOUT_TEMPR79[6] , 
        \B_DOUT_TEMPR80[6] , \B_DOUT_TEMPR81[6] , \B_DOUT_TEMPR82[6] , 
        \B_DOUT_TEMPR83[6] , \B_DOUT_TEMPR84[6] , \B_DOUT_TEMPR85[6] , 
        \B_DOUT_TEMPR86[6] , \B_DOUT_TEMPR87[6] , \B_DOUT_TEMPR88[6] , 
        \B_DOUT_TEMPR89[6] , \B_DOUT_TEMPR90[6] , \B_DOUT_TEMPR91[6] , 
        \B_DOUT_TEMPR92[6] , \B_DOUT_TEMPR93[6] , \B_DOUT_TEMPR94[6] , 
        \B_DOUT_TEMPR95[6] , \B_DOUT_TEMPR96[6] , \B_DOUT_TEMPR97[6] , 
        \B_DOUT_TEMPR98[6] , \B_DOUT_TEMPR99[6] , \B_DOUT_TEMPR100[6] , 
        \B_DOUT_TEMPR101[6] , \B_DOUT_TEMPR102[6] , 
        \B_DOUT_TEMPR103[6] , \B_DOUT_TEMPR104[6] , 
        \B_DOUT_TEMPR105[6] , \B_DOUT_TEMPR106[6] , 
        \B_DOUT_TEMPR107[6] , \B_DOUT_TEMPR108[6] , 
        \B_DOUT_TEMPR109[6] , \B_DOUT_TEMPR110[6] , 
        \B_DOUT_TEMPR111[6] , \B_DOUT_TEMPR112[6] , 
        \B_DOUT_TEMPR113[6] , \B_DOUT_TEMPR114[6] , 
        \B_DOUT_TEMPR115[6] , \B_DOUT_TEMPR116[6] , 
        \B_DOUT_TEMPR117[6] , \B_DOUT_TEMPR118[6] , \B_DOUT_TEMPR0[7] , 
        \B_DOUT_TEMPR1[7] , \B_DOUT_TEMPR2[7] , \B_DOUT_TEMPR3[7] , 
        \B_DOUT_TEMPR4[7] , \B_DOUT_TEMPR5[7] , \B_DOUT_TEMPR6[7] , 
        \B_DOUT_TEMPR7[7] , \B_DOUT_TEMPR8[7] , \B_DOUT_TEMPR9[7] , 
        \B_DOUT_TEMPR10[7] , \B_DOUT_TEMPR11[7] , \B_DOUT_TEMPR12[7] , 
        \B_DOUT_TEMPR13[7] , \B_DOUT_TEMPR14[7] , \B_DOUT_TEMPR15[7] , 
        \B_DOUT_TEMPR16[7] , \B_DOUT_TEMPR17[7] , \B_DOUT_TEMPR18[7] , 
        \B_DOUT_TEMPR19[7] , \B_DOUT_TEMPR20[7] , \B_DOUT_TEMPR21[7] , 
        \B_DOUT_TEMPR22[7] , \B_DOUT_TEMPR23[7] , \B_DOUT_TEMPR24[7] , 
        \B_DOUT_TEMPR25[7] , \B_DOUT_TEMPR26[7] , \B_DOUT_TEMPR27[7] , 
        \B_DOUT_TEMPR28[7] , \B_DOUT_TEMPR29[7] , \B_DOUT_TEMPR30[7] , 
        \B_DOUT_TEMPR31[7] , \B_DOUT_TEMPR32[7] , \B_DOUT_TEMPR33[7] , 
        \B_DOUT_TEMPR34[7] , \B_DOUT_TEMPR35[7] , \B_DOUT_TEMPR36[7] , 
        \B_DOUT_TEMPR37[7] , \B_DOUT_TEMPR38[7] , \B_DOUT_TEMPR39[7] , 
        \B_DOUT_TEMPR40[7] , \B_DOUT_TEMPR41[7] , \B_DOUT_TEMPR42[7] , 
        \B_DOUT_TEMPR43[7] , \B_DOUT_TEMPR44[7] , \B_DOUT_TEMPR45[7] , 
        \B_DOUT_TEMPR46[7] , \B_DOUT_TEMPR47[7] , \B_DOUT_TEMPR48[7] , 
        \B_DOUT_TEMPR49[7] , \B_DOUT_TEMPR50[7] , \B_DOUT_TEMPR51[7] , 
        \B_DOUT_TEMPR52[7] , \B_DOUT_TEMPR53[7] , \B_DOUT_TEMPR54[7] , 
        \B_DOUT_TEMPR55[7] , \B_DOUT_TEMPR56[7] , \B_DOUT_TEMPR57[7] , 
        \B_DOUT_TEMPR58[7] , \B_DOUT_TEMPR59[7] , \B_DOUT_TEMPR60[7] , 
        \B_DOUT_TEMPR61[7] , \B_DOUT_TEMPR62[7] , \B_DOUT_TEMPR63[7] , 
        \B_DOUT_TEMPR64[7] , \B_DOUT_TEMPR65[7] , \B_DOUT_TEMPR66[7] , 
        \B_DOUT_TEMPR67[7] , \B_DOUT_TEMPR68[7] , \B_DOUT_TEMPR69[7] , 
        \B_DOUT_TEMPR70[7] , \B_DOUT_TEMPR71[7] , \B_DOUT_TEMPR72[7] , 
        \B_DOUT_TEMPR73[7] , \B_DOUT_TEMPR74[7] , \B_DOUT_TEMPR75[7] , 
        \B_DOUT_TEMPR76[7] , \B_DOUT_TEMPR77[7] , \B_DOUT_TEMPR78[7] , 
        \B_DOUT_TEMPR79[7] , \B_DOUT_TEMPR80[7] , \B_DOUT_TEMPR81[7] , 
        \B_DOUT_TEMPR82[7] , \B_DOUT_TEMPR83[7] , \B_DOUT_TEMPR84[7] , 
        \B_DOUT_TEMPR85[7] , \B_DOUT_TEMPR86[7] , \B_DOUT_TEMPR87[7] , 
        \B_DOUT_TEMPR88[7] , \B_DOUT_TEMPR89[7] , \B_DOUT_TEMPR90[7] , 
        \B_DOUT_TEMPR91[7] , \B_DOUT_TEMPR92[7] , \B_DOUT_TEMPR93[7] , 
        \B_DOUT_TEMPR94[7] , \B_DOUT_TEMPR95[7] , \B_DOUT_TEMPR96[7] , 
        \B_DOUT_TEMPR97[7] , \B_DOUT_TEMPR98[7] , \B_DOUT_TEMPR99[7] , 
        \B_DOUT_TEMPR100[7] , \B_DOUT_TEMPR101[7] , 
        \B_DOUT_TEMPR102[7] , \B_DOUT_TEMPR103[7] , 
        \B_DOUT_TEMPR104[7] , \B_DOUT_TEMPR105[7] , 
        \B_DOUT_TEMPR106[7] , \B_DOUT_TEMPR107[7] , 
        \B_DOUT_TEMPR108[7] , \B_DOUT_TEMPR109[7] , 
        \B_DOUT_TEMPR110[7] , \B_DOUT_TEMPR111[7] , 
        \B_DOUT_TEMPR112[7] , \B_DOUT_TEMPR113[7] , 
        \B_DOUT_TEMPR114[7] , \B_DOUT_TEMPR115[7] , 
        \B_DOUT_TEMPR116[7] , \B_DOUT_TEMPR117[7] , 
        \B_DOUT_TEMPR118[7] , \B_DOUT_TEMPR0[8] , \B_DOUT_TEMPR1[8] , 
        \B_DOUT_TEMPR2[8] , \B_DOUT_TEMPR3[8] , \B_DOUT_TEMPR4[8] , 
        \B_DOUT_TEMPR5[8] , \B_DOUT_TEMPR6[8] , \B_DOUT_TEMPR7[8] , 
        \B_DOUT_TEMPR8[8] , \B_DOUT_TEMPR9[8] , \B_DOUT_TEMPR10[8] , 
        \B_DOUT_TEMPR11[8] , \B_DOUT_TEMPR12[8] , \B_DOUT_TEMPR13[8] , 
        \B_DOUT_TEMPR14[8] , \B_DOUT_TEMPR15[8] , \B_DOUT_TEMPR16[8] , 
        \B_DOUT_TEMPR17[8] , \B_DOUT_TEMPR18[8] , \B_DOUT_TEMPR19[8] , 
        \B_DOUT_TEMPR20[8] , \B_DOUT_TEMPR21[8] , \B_DOUT_TEMPR22[8] , 
        \B_DOUT_TEMPR23[8] , \B_DOUT_TEMPR24[8] , \B_DOUT_TEMPR25[8] , 
        \B_DOUT_TEMPR26[8] , \B_DOUT_TEMPR27[8] , \B_DOUT_TEMPR28[8] , 
        \B_DOUT_TEMPR29[8] , \B_DOUT_TEMPR30[8] , \B_DOUT_TEMPR31[8] , 
        \B_DOUT_TEMPR32[8] , \B_DOUT_TEMPR33[8] , \B_DOUT_TEMPR34[8] , 
        \B_DOUT_TEMPR35[8] , \B_DOUT_TEMPR36[8] , \B_DOUT_TEMPR37[8] , 
        \B_DOUT_TEMPR38[8] , \B_DOUT_TEMPR39[8] , \B_DOUT_TEMPR40[8] , 
        \B_DOUT_TEMPR41[8] , \B_DOUT_TEMPR42[8] , \B_DOUT_TEMPR43[8] , 
        \B_DOUT_TEMPR44[8] , \B_DOUT_TEMPR45[8] , \B_DOUT_TEMPR46[8] , 
        \B_DOUT_TEMPR47[8] , \B_DOUT_TEMPR48[8] , \B_DOUT_TEMPR49[8] , 
        \B_DOUT_TEMPR50[8] , \B_DOUT_TEMPR51[8] , \B_DOUT_TEMPR52[8] , 
        \B_DOUT_TEMPR53[8] , \B_DOUT_TEMPR54[8] , \B_DOUT_TEMPR55[8] , 
        \B_DOUT_TEMPR56[8] , \B_DOUT_TEMPR57[8] , \B_DOUT_TEMPR58[8] , 
        \B_DOUT_TEMPR59[8] , \B_DOUT_TEMPR60[8] , \B_DOUT_TEMPR61[8] , 
        \B_DOUT_TEMPR62[8] , \B_DOUT_TEMPR63[8] , \B_DOUT_TEMPR64[8] , 
        \B_DOUT_TEMPR65[8] , \B_DOUT_TEMPR66[8] , \B_DOUT_TEMPR67[8] , 
        \B_DOUT_TEMPR68[8] , \B_DOUT_TEMPR69[8] , \B_DOUT_TEMPR70[8] , 
        \B_DOUT_TEMPR71[8] , \B_DOUT_TEMPR72[8] , \B_DOUT_TEMPR73[8] , 
        \B_DOUT_TEMPR74[8] , \B_DOUT_TEMPR75[8] , \B_DOUT_TEMPR76[8] , 
        \B_DOUT_TEMPR77[8] , \B_DOUT_TEMPR78[8] , \B_DOUT_TEMPR79[8] , 
        \B_DOUT_TEMPR80[8] , \B_DOUT_TEMPR81[8] , \B_DOUT_TEMPR82[8] , 
        \B_DOUT_TEMPR83[8] , \B_DOUT_TEMPR84[8] , \B_DOUT_TEMPR85[8] , 
        \B_DOUT_TEMPR86[8] , \B_DOUT_TEMPR87[8] , \B_DOUT_TEMPR88[8] , 
        \B_DOUT_TEMPR89[8] , \B_DOUT_TEMPR90[8] , \B_DOUT_TEMPR91[8] , 
        \B_DOUT_TEMPR92[8] , \B_DOUT_TEMPR93[8] , \B_DOUT_TEMPR94[8] , 
        \B_DOUT_TEMPR95[8] , \B_DOUT_TEMPR96[8] , \B_DOUT_TEMPR97[8] , 
        \B_DOUT_TEMPR98[8] , \B_DOUT_TEMPR99[8] , \B_DOUT_TEMPR100[8] , 
        \B_DOUT_TEMPR101[8] , \B_DOUT_TEMPR102[8] , 
        \B_DOUT_TEMPR103[8] , \B_DOUT_TEMPR104[8] , 
        \B_DOUT_TEMPR105[8] , \B_DOUT_TEMPR106[8] , 
        \B_DOUT_TEMPR107[8] , \B_DOUT_TEMPR108[8] , 
        \B_DOUT_TEMPR109[8] , \B_DOUT_TEMPR110[8] , 
        \B_DOUT_TEMPR111[8] , \B_DOUT_TEMPR112[8] , 
        \B_DOUT_TEMPR113[8] , \B_DOUT_TEMPR114[8] , 
        \B_DOUT_TEMPR115[8] , \B_DOUT_TEMPR116[8] , 
        \B_DOUT_TEMPR117[8] , \B_DOUT_TEMPR118[8] , \B_DOUT_TEMPR0[9] , 
        \B_DOUT_TEMPR1[9] , \B_DOUT_TEMPR2[9] , \B_DOUT_TEMPR3[9] , 
        \B_DOUT_TEMPR4[9] , \B_DOUT_TEMPR5[9] , \B_DOUT_TEMPR6[9] , 
        \B_DOUT_TEMPR7[9] , \B_DOUT_TEMPR8[9] , \B_DOUT_TEMPR9[9] , 
        \B_DOUT_TEMPR10[9] , \B_DOUT_TEMPR11[9] , \B_DOUT_TEMPR12[9] , 
        \B_DOUT_TEMPR13[9] , \B_DOUT_TEMPR14[9] , \B_DOUT_TEMPR15[9] , 
        \B_DOUT_TEMPR16[9] , \B_DOUT_TEMPR17[9] , \B_DOUT_TEMPR18[9] , 
        \B_DOUT_TEMPR19[9] , \B_DOUT_TEMPR20[9] , \B_DOUT_TEMPR21[9] , 
        \B_DOUT_TEMPR22[9] , \B_DOUT_TEMPR23[9] , \B_DOUT_TEMPR24[9] , 
        \B_DOUT_TEMPR25[9] , \B_DOUT_TEMPR26[9] , \B_DOUT_TEMPR27[9] , 
        \B_DOUT_TEMPR28[9] , \B_DOUT_TEMPR29[9] , \B_DOUT_TEMPR30[9] , 
        \B_DOUT_TEMPR31[9] , \B_DOUT_TEMPR32[9] , \B_DOUT_TEMPR33[9] , 
        \B_DOUT_TEMPR34[9] , \B_DOUT_TEMPR35[9] , \B_DOUT_TEMPR36[9] , 
        \B_DOUT_TEMPR37[9] , \B_DOUT_TEMPR38[9] , \B_DOUT_TEMPR39[9] , 
        \B_DOUT_TEMPR40[9] , \B_DOUT_TEMPR41[9] , \B_DOUT_TEMPR42[9] , 
        \B_DOUT_TEMPR43[9] , \B_DOUT_TEMPR44[9] , \B_DOUT_TEMPR45[9] , 
        \B_DOUT_TEMPR46[9] , \B_DOUT_TEMPR47[9] , \B_DOUT_TEMPR48[9] , 
        \B_DOUT_TEMPR49[9] , \B_DOUT_TEMPR50[9] , \B_DOUT_TEMPR51[9] , 
        \B_DOUT_TEMPR52[9] , \B_DOUT_TEMPR53[9] , \B_DOUT_TEMPR54[9] , 
        \B_DOUT_TEMPR55[9] , \B_DOUT_TEMPR56[9] , \B_DOUT_TEMPR57[9] , 
        \B_DOUT_TEMPR58[9] , \B_DOUT_TEMPR59[9] , \B_DOUT_TEMPR60[9] , 
        \B_DOUT_TEMPR61[9] , \B_DOUT_TEMPR62[9] , \B_DOUT_TEMPR63[9] , 
        \B_DOUT_TEMPR64[9] , \B_DOUT_TEMPR65[9] , \B_DOUT_TEMPR66[9] , 
        \B_DOUT_TEMPR67[9] , \B_DOUT_TEMPR68[9] , \B_DOUT_TEMPR69[9] , 
        \B_DOUT_TEMPR70[9] , \B_DOUT_TEMPR71[9] , \B_DOUT_TEMPR72[9] , 
        \B_DOUT_TEMPR73[9] , \B_DOUT_TEMPR74[9] , \B_DOUT_TEMPR75[9] , 
        \B_DOUT_TEMPR76[9] , \B_DOUT_TEMPR77[9] , \B_DOUT_TEMPR78[9] , 
        \B_DOUT_TEMPR79[9] , \B_DOUT_TEMPR80[9] , \B_DOUT_TEMPR81[9] , 
        \B_DOUT_TEMPR82[9] , \B_DOUT_TEMPR83[9] , \B_DOUT_TEMPR84[9] , 
        \B_DOUT_TEMPR85[9] , \B_DOUT_TEMPR86[9] , \B_DOUT_TEMPR87[9] , 
        \B_DOUT_TEMPR88[9] , \B_DOUT_TEMPR89[9] , \B_DOUT_TEMPR90[9] , 
        \B_DOUT_TEMPR91[9] , \B_DOUT_TEMPR92[9] , \B_DOUT_TEMPR93[9] , 
        \B_DOUT_TEMPR94[9] , \B_DOUT_TEMPR95[9] , \B_DOUT_TEMPR96[9] , 
        \B_DOUT_TEMPR97[9] , \B_DOUT_TEMPR98[9] , \B_DOUT_TEMPR99[9] , 
        \B_DOUT_TEMPR100[9] , \B_DOUT_TEMPR101[9] , 
        \B_DOUT_TEMPR102[9] , \B_DOUT_TEMPR103[9] , 
        \B_DOUT_TEMPR104[9] , \B_DOUT_TEMPR105[9] , 
        \B_DOUT_TEMPR106[9] , \B_DOUT_TEMPR107[9] , 
        \B_DOUT_TEMPR108[9] , \B_DOUT_TEMPR109[9] , 
        \B_DOUT_TEMPR110[9] , \B_DOUT_TEMPR111[9] , 
        \B_DOUT_TEMPR112[9] , \B_DOUT_TEMPR113[9] , 
        \B_DOUT_TEMPR114[9] , \B_DOUT_TEMPR115[9] , 
        \B_DOUT_TEMPR116[9] , \B_DOUT_TEMPR117[9] , 
        \B_DOUT_TEMPR118[9] , \B_DOUT_TEMPR0[10] , \B_DOUT_TEMPR1[10] , 
        \B_DOUT_TEMPR2[10] , \B_DOUT_TEMPR3[10] , \B_DOUT_TEMPR4[10] , 
        \B_DOUT_TEMPR5[10] , \B_DOUT_TEMPR6[10] , \B_DOUT_TEMPR7[10] , 
        \B_DOUT_TEMPR8[10] , \B_DOUT_TEMPR9[10] , \B_DOUT_TEMPR10[10] , 
        \B_DOUT_TEMPR11[10] , \B_DOUT_TEMPR12[10] , 
        \B_DOUT_TEMPR13[10] , \B_DOUT_TEMPR14[10] , 
        \B_DOUT_TEMPR15[10] , \B_DOUT_TEMPR16[10] , 
        \B_DOUT_TEMPR17[10] , \B_DOUT_TEMPR18[10] , 
        \B_DOUT_TEMPR19[10] , \B_DOUT_TEMPR20[10] , 
        \B_DOUT_TEMPR21[10] , \B_DOUT_TEMPR22[10] , 
        \B_DOUT_TEMPR23[10] , \B_DOUT_TEMPR24[10] , 
        \B_DOUT_TEMPR25[10] , \B_DOUT_TEMPR26[10] , 
        \B_DOUT_TEMPR27[10] , \B_DOUT_TEMPR28[10] , 
        \B_DOUT_TEMPR29[10] , \B_DOUT_TEMPR30[10] , 
        \B_DOUT_TEMPR31[10] , \B_DOUT_TEMPR32[10] , 
        \B_DOUT_TEMPR33[10] , \B_DOUT_TEMPR34[10] , 
        \B_DOUT_TEMPR35[10] , \B_DOUT_TEMPR36[10] , 
        \B_DOUT_TEMPR37[10] , \B_DOUT_TEMPR38[10] , 
        \B_DOUT_TEMPR39[10] , \B_DOUT_TEMPR40[10] , 
        \B_DOUT_TEMPR41[10] , \B_DOUT_TEMPR42[10] , 
        \B_DOUT_TEMPR43[10] , \B_DOUT_TEMPR44[10] , 
        \B_DOUT_TEMPR45[10] , \B_DOUT_TEMPR46[10] , 
        \B_DOUT_TEMPR47[10] , \B_DOUT_TEMPR48[10] , 
        \B_DOUT_TEMPR49[10] , \B_DOUT_TEMPR50[10] , 
        \B_DOUT_TEMPR51[10] , \B_DOUT_TEMPR52[10] , 
        \B_DOUT_TEMPR53[10] , \B_DOUT_TEMPR54[10] , 
        \B_DOUT_TEMPR55[10] , \B_DOUT_TEMPR56[10] , 
        \B_DOUT_TEMPR57[10] , \B_DOUT_TEMPR58[10] , 
        \B_DOUT_TEMPR59[10] , \B_DOUT_TEMPR60[10] , 
        \B_DOUT_TEMPR61[10] , \B_DOUT_TEMPR62[10] , 
        \B_DOUT_TEMPR63[10] , \B_DOUT_TEMPR64[10] , 
        \B_DOUT_TEMPR65[10] , \B_DOUT_TEMPR66[10] , 
        \B_DOUT_TEMPR67[10] , \B_DOUT_TEMPR68[10] , 
        \B_DOUT_TEMPR69[10] , \B_DOUT_TEMPR70[10] , 
        \B_DOUT_TEMPR71[10] , \B_DOUT_TEMPR72[10] , 
        \B_DOUT_TEMPR73[10] , \B_DOUT_TEMPR74[10] , 
        \B_DOUT_TEMPR75[10] , \B_DOUT_TEMPR76[10] , 
        \B_DOUT_TEMPR77[10] , \B_DOUT_TEMPR78[10] , 
        \B_DOUT_TEMPR79[10] , \B_DOUT_TEMPR80[10] , 
        \B_DOUT_TEMPR81[10] , \B_DOUT_TEMPR82[10] , 
        \B_DOUT_TEMPR83[10] , \B_DOUT_TEMPR84[10] , 
        \B_DOUT_TEMPR85[10] , \B_DOUT_TEMPR86[10] , 
        \B_DOUT_TEMPR87[10] , \B_DOUT_TEMPR88[10] , 
        \B_DOUT_TEMPR89[10] , \B_DOUT_TEMPR90[10] , 
        \B_DOUT_TEMPR91[10] , \B_DOUT_TEMPR92[10] , 
        \B_DOUT_TEMPR93[10] , \B_DOUT_TEMPR94[10] , 
        \B_DOUT_TEMPR95[10] , \B_DOUT_TEMPR96[10] , 
        \B_DOUT_TEMPR97[10] , \B_DOUT_TEMPR98[10] , 
        \B_DOUT_TEMPR99[10] , \B_DOUT_TEMPR100[10] , 
        \B_DOUT_TEMPR101[10] , \B_DOUT_TEMPR102[10] , 
        \B_DOUT_TEMPR103[10] , \B_DOUT_TEMPR104[10] , 
        \B_DOUT_TEMPR105[10] , \B_DOUT_TEMPR106[10] , 
        \B_DOUT_TEMPR107[10] , \B_DOUT_TEMPR108[10] , 
        \B_DOUT_TEMPR109[10] , \B_DOUT_TEMPR110[10] , 
        \B_DOUT_TEMPR111[10] , \B_DOUT_TEMPR112[10] , 
        \B_DOUT_TEMPR113[10] , \B_DOUT_TEMPR114[10] , 
        \B_DOUT_TEMPR115[10] , \B_DOUT_TEMPR116[10] , 
        \B_DOUT_TEMPR117[10] , \B_DOUT_TEMPR118[10] , 
        \B_DOUT_TEMPR0[11] , \B_DOUT_TEMPR1[11] , \B_DOUT_TEMPR2[11] , 
        \B_DOUT_TEMPR3[11] , \B_DOUT_TEMPR4[11] , \B_DOUT_TEMPR5[11] , 
        \B_DOUT_TEMPR6[11] , \B_DOUT_TEMPR7[11] , \B_DOUT_TEMPR8[11] , 
        \B_DOUT_TEMPR9[11] , \B_DOUT_TEMPR10[11] , 
        \B_DOUT_TEMPR11[11] , \B_DOUT_TEMPR12[11] , 
        \B_DOUT_TEMPR13[11] , \B_DOUT_TEMPR14[11] , 
        \B_DOUT_TEMPR15[11] , \B_DOUT_TEMPR16[11] , 
        \B_DOUT_TEMPR17[11] , \B_DOUT_TEMPR18[11] , 
        \B_DOUT_TEMPR19[11] , \B_DOUT_TEMPR20[11] , 
        \B_DOUT_TEMPR21[11] , \B_DOUT_TEMPR22[11] , 
        \B_DOUT_TEMPR23[11] , \B_DOUT_TEMPR24[11] , 
        \B_DOUT_TEMPR25[11] , \B_DOUT_TEMPR26[11] , 
        \B_DOUT_TEMPR27[11] , \B_DOUT_TEMPR28[11] , 
        \B_DOUT_TEMPR29[11] , \B_DOUT_TEMPR30[11] , 
        \B_DOUT_TEMPR31[11] , \B_DOUT_TEMPR32[11] , 
        \B_DOUT_TEMPR33[11] , \B_DOUT_TEMPR34[11] , 
        \B_DOUT_TEMPR35[11] , \B_DOUT_TEMPR36[11] , 
        \B_DOUT_TEMPR37[11] , \B_DOUT_TEMPR38[11] , 
        \B_DOUT_TEMPR39[11] , \B_DOUT_TEMPR40[11] , 
        \B_DOUT_TEMPR41[11] , \B_DOUT_TEMPR42[11] , 
        \B_DOUT_TEMPR43[11] , \B_DOUT_TEMPR44[11] , 
        \B_DOUT_TEMPR45[11] , \B_DOUT_TEMPR46[11] , 
        \B_DOUT_TEMPR47[11] , \B_DOUT_TEMPR48[11] , 
        \B_DOUT_TEMPR49[11] , \B_DOUT_TEMPR50[11] , 
        \B_DOUT_TEMPR51[11] , \B_DOUT_TEMPR52[11] , 
        \B_DOUT_TEMPR53[11] , \B_DOUT_TEMPR54[11] , 
        \B_DOUT_TEMPR55[11] , \B_DOUT_TEMPR56[11] , 
        \B_DOUT_TEMPR57[11] , \B_DOUT_TEMPR58[11] , 
        \B_DOUT_TEMPR59[11] , \B_DOUT_TEMPR60[11] , 
        \B_DOUT_TEMPR61[11] , \B_DOUT_TEMPR62[11] , 
        \B_DOUT_TEMPR63[11] , \B_DOUT_TEMPR64[11] , 
        \B_DOUT_TEMPR65[11] , \B_DOUT_TEMPR66[11] , 
        \B_DOUT_TEMPR67[11] , \B_DOUT_TEMPR68[11] , 
        \B_DOUT_TEMPR69[11] , \B_DOUT_TEMPR70[11] , 
        \B_DOUT_TEMPR71[11] , \B_DOUT_TEMPR72[11] , 
        \B_DOUT_TEMPR73[11] , \B_DOUT_TEMPR74[11] , 
        \B_DOUT_TEMPR75[11] , \B_DOUT_TEMPR76[11] , 
        \B_DOUT_TEMPR77[11] , \B_DOUT_TEMPR78[11] , 
        \B_DOUT_TEMPR79[11] , \B_DOUT_TEMPR80[11] , 
        \B_DOUT_TEMPR81[11] , \B_DOUT_TEMPR82[11] , 
        \B_DOUT_TEMPR83[11] , \B_DOUT_TEMPR84[11] , 
        \B_DOUT_TEMPR85[11] , \B_DOUT_TEMPR86[11] , 
        \B_DOUT_TEMPR87[11] , \B_DOUT_TEMPR88[11] , 
        \B_DOUT_TEMPR89[11] , \B_DOUT_TEMPR90[11] , 
        \B_DOUT_TEMPR91[11] , \B_DOUT_TEMPR92[11] , 
        \B_DOUT_TEMPR93[11] , \B_DOUT_TEMPR94[11] , 
        \B_DOUT_TEMPR95[11] , \B_DOUT_TEMPR96[11] , 
        \B_DOUT_TEMPR97[11] , \B_DOUT_TEMPR98[11] , 
        \B_DOUT_TEMPR99[11] , \B_DOUT_TEMPR100[11] , 
        \B_DOUT_TEMPR101[11] , \B_DOUT_TEMPR102[11] , 
        \B_DOUT_TEMPR103[11] , \B_DOUT_TEMPR104[11] , 
        \B_DOUT_TEMPR105[11] , \B_DOUT_TEMPR106[11] , 
        \B_DOUT_TEMPR107[11] , \B_DOUT_TEMPR108[11] , 
        \B_DOUT_TEMPR109[11] , \B_DOUT_TEMPR110[11] , 
        \B_DOUT_TEMPR111[11] , \B_DOUT_TEMPR112[11] , 
        \B_DOUT_TEMPR113[11] , \B_DOUT_TEMPR114[11] , 
        \B_DOUT_TEMPR115[11] , \B_DOUT_TEMPR116[11] , 
        \B_DOUT_TEMPR117[11] , \B_DOUT_TEMPR118[11] , 
        \B_DOUT_TEMPR0[12] , \B_DOUT_TEMPR1[12] , \B_DOUT_TEMPR2[12] , 
        \B_DOUT_TEMPR3[12] , \B_DOUT_TEMPR4[12] , \B_DOUT_TEMPR5[12] , 
        \B_DOUT_TEMPR6[12] , \B_DOUT_TEMPR7[12] , \B_DOUT_TEMPR8[12] , 
        \B_DOUT_TEMPR9[12] , \B_DOUT_TEMPR10[12] , 
        \B_DOUT_TEMPR11[12] , \B_DOUT_TEMPR12[12] , 
        \B_DOUT_TEMPR13[12] , \B_DOUT_TEMPR14[12] , 
        \B_DOUT_TEMPR15[12] , \B_DOUT_TEMPR16[12] , 
        \B_DOUT_TEMPR17[12] , \B_DOUT_TEMPR18[12] , 
        \B_DOUT_TEMPR19[12] , \B_DOUT_TEMPR20[12] , 
        \B_DOUT_TEMPR21[12] , \B_DOUT_TEMPR22[12] , 
        \B_DOUT_TEMPR23[12] , \B_DOUT_TEMPR24[12] , 
        \B_DOUT_TEMPR25[12] , \B_DOUT_TEMPR26[12] , 
        \B_DOUT_TEMPR27[12] , \B_DOUT_TEMPR28[12] , 
        \B_DOUT_TEMPR29[12] , \B_DOUT_TEMPR30[12] , 
        \B_DOUT_TEMPR31[12] , \B_DOUT_TEMPR32[12] , 
        \B_DOUT_TEMPR33[12] , \B_DOUT_TEMPR34[12] , 
        \B_DOUT_TEMPR35[12] , \B_DOUT_TEMPR36[12] , 
        \B_DOUT_TEMPR37[12] , \B_DOUT_TEMPR38[12] , 
        \B_DOUT_TEMPR39[12] , \B_DOUT_TEMPR40[12] , 
        \B_DOUT_TEMPR41[12] , \B_DOUT_TEMPR42[12] , 
        \B_DOUT_TEMPR43[12] , \B_DOUT_TEMPR44[12] , 
        \B_DOUT_TEMPR45[12] , \B_DOUT_TEMPR46[12] , 
        \B_DOUT_TEMPR47[12] , \B_DOUT_TEMPR48[12] , 
        \B_DOUT_TEMPR49[12] , \B_DOUT_TEMPR50[12] , 
        \B_DOUT_TEMPR51[12] , \B_DOUT_TEMPR52[12] , 
        \B_DOUT_TEMPR53[12] , \B_DOUT_TEMPR54[12] , 
        \B_DOUT_TEMPR55[12] , \B_DOUT_TEMPR56[12] , 
        \B_DOUT_TEMPR57[12] , \B_DOUT_TEMPR58[12] , 
        \B_DOUT_TEMPR59[12] , \B_DOUT_TEMPR60[12] , 
        \B_DOUT_TEMPR61[12] , \B_DOUT_TEMPR62[12] , 
        \B_DOUT_TEMPR63[12] , \B_DOUT_TEMPR64[12] , 
        \B_DOUT_TEMPR65[12] , \B_DOUT_TEMPR66[12] , 
        \B_DOUT_TEMPR67[12] , \B_DOUT_TEMPR68[12] , 
        \B_DOUT_TEMPR69[12] , \B_DOUT_TEMPR70[12] , 
        \B_DOUT_TEMPR71[12] , \B_DOUT_TEMPR72[12] , 
        \B_DOUT_TEMPR73[12] , \B_DOUT_TEMPR74[12] , 
        \B_DOUT_TEMPR75[12] , \B_DOUT_TEMPR76[12] , 
        \B_DOUT_TEMPR77[12] , \B_DOUT_TEMPR78[12] , 
        \B_DOUT_TEMPR79[12] , \B_DOUT_TEMPR80[12] , 
        \B_DOUT_TEMPR81[12] , \B_DOUT_TEMPR82[12] , 
        \B_DOUT_TEMPR83[12] , \B_DOUT_TEMPR84[12] , 
        \B_DOUT_TEMPR85[12] , \B_DOUT_TEMPR86[12] , 
        \B_DOUT_TEMPR87[12] , \B_DOUT_TEMPR88[12] , 
        \B_DOUT_TEMPR89[12] , \B_DOUT_TEMPR90[12] , 
        \B_DOUT_TEMPR91[12] , \B_DOUT_TEMPR92[12] , 
        \B_DOUT_TEMPR93[12] , \B_DOUT_TEMPR94[12] , 
        \B_DOUT_TEMPR95[12] , \B_DOUT_TEMPR96[12] , 
        \B_DOUT_TEMPR97[12] , \B_DOUT_TEMPR98[12] , 
        \B_DOUT_TEMPR99[12] , \B_DOUT_TEMPR100[12] , 
        \B_DOUT_TEMPR101[12] , \B_DOUT_TEMPR102[12] , 
        \B_DOUT_TEMPR103[12] , \B_DOUT_TEMPR104[12] , 
        \B_DOUT_TEMPR105[12] , \B_DOUT_TEMPR106[12] , 
        \B_DOUT_TEMPR107[12] , \B_DOUT_TEMPR108[12] , 
        \B_DOUT_TEMPR109[12] , \B_DOUT_TEMPR110[12] , 
        \B_DOUT_TEMPR111[12] , \B_DOUT_TEMPR112[12] , 
        \B_DOUT_TEMPR113[12] , \B_DOUT_TEMPR114[12] , 
        \B_DOUT_TEMPR115[12] , \B_DOUT_TEMPR116[12] , 
        \B_DOUT_TEMPR117[12] , \B_DOUT_TEMPR118[12] , 
        \B_DOUT_TEMPR0[13] , \B_DOUT_TEMPR1[13] , \B_DOUT_TEMPR2[13] , 
        \B_DOUT_TEMPR3[13] , \B_DOUT_TEMPR4[13] , \B_DOUT_TEMPR5[13] , 
        \B_DOUT_TEMPR6[13] , \B_DOUT_TEMPR7[13] , \B_DOUT_TEMPR8[13] , 
        \B_DOUT_TEMPR9[13] , \B_DOUT_TEMPR10[13] , 
        \B_DOUT_TEMPR11[13] , \B_DOUT_TEMPR12[13] , 
        \B_DOUT_TEMPR13[13] , \B_DOUT_TEMPR14[13] , 
        \B_DOUT_TEMPR15[13] , \B_DOUT_TEMPR16[13] , 
        \B_DOUT_TEMPR17[13] , \B_DOUT_TEMPR18[13] , 
        \B_DOUT_TEMPR19[13] , \B_DOUT_TEMPR20[13] , 
        \B_DOUT_TEMPR21[13] , \B_DOUT_TEMPR22[13] , 
        \B_DOUT_TEMPR23[13] , \B_DOUT_TEMPR24[13] , 
        \B_DOUT_TEMPR25[13] , \B_DOUT_TEMPR26[13] , 
        \B_DOUT_TEMPR27[13] , \B_DOUT_TEMPR28[13] , 
        \B_DOUT_TEMPR29[13] , \B_DOUT_TEMPR30[13] , 
        \B_DOUT_TEMPR31[13] , \B_DOUT_TEMPR32[13] , 
        \B_DOUT_TEMPR33[13] , \B_DOUT_TEMPR34[13] , 
        \B_DOUT_TEMPR35[13] , \B_DOUT_TEMPR36[13] , 
        \B_DOUT_TEMPR37[13] , \B_DOUT_TEMPR38[13] , 
        \B_DOUT_TEMPR39[13] , \B_DOUT_TEMPR40[13] , 
        \B_DOUT_TEMPR41[13] , \B_DOUT_TEMPR42[13] , 
        \B_DOUT_TEMPR43[13] , \B_DOUT_TEMPR44[13] , 
        \B_DOUT_TEMPR45[13] , \B_DOUT_TEMPR46[13] , 
        \B_DOUT_TEMPR47[13] , \B_DOUT_TEMPR48[13] , 
        \B_DOUT_TEMPR49[13] , \B_DOUT_TEMPR50[13] , 
        \B_DOUT_TEMPR51[13] , \B_DOUT_TEMPR52[13] , 
        \B_DOUT_TEMPR53[13] , \B_DOUT_TEMPR54[13] , 
        \B_DOUT_TEMPR55[13] , \B_DOUT_TEMPR56[13] , 
        \B_DOUT_TEMPR57[13] , \B_DOUT_TEMPR58[13] , 
        \B_DOUT_TEMPR59[13] , \B_DOUT_TEMPR60[13] , 
        \B_DOUT_TEMPR61[13] , \B_DOUT_TEMPR62[13] , 
        \B_DOUT_TEMPR63[13] , \B_DOUT_TEMPR64[13] , 
        \B_DOUT_TEMPR65[13] , \B_DOUT_TEMPR66[13] , 
        \B_DOUT_TEMPR67[13] , \B_DOUT_TEMPR68[13] , 
        \B_DOUT_TEMPR69[13] , \B_DOUT_TEMPR70[13] , 
        \B_DOUT_TEMPR71[13] , \B_DOUT_TEMPR72[13] , 
        \B_DOUT_TEMPR73[13] , \B_DOUT_TEMPR74[13] , 
        \B_DOUT_TEMPR75[13] , \B_DOUT_TEMPR76[13] , 
        \B_DOUT_TEMPR77[13] , \B_DOUT_TEMPR78[13] , 
        \B_DOUT_TEMPR79[13] , \B_DOUT_TEMPR80[13] , 
        \B_DOUT_TEMPR81[13] , \B_DOUT_TEMPR82[13] , 
        \B_DOUT_TEMPR83[13] , \B_DOUT_TEMPR84[13] , 
        \B_DOUT_TEMPR85[13] , \B_DOUT_TEMPR86[13] , 
        \B_DOUT_TEMPR87[13] , \B_DOUT_TEMPR88[13] , 
        \B_DOUT_TEMPR89[13] , \B_DOUT_TEMPR90[13] , 
        \B_DOUT_TEMPR91[13] , \B_DOUT_TEMPR92[13] , 
        \B_DOUT_TEMPR93[13] , \B_DOUT_TEMPR94[13] , 
        \B_DOUT_TEMPR95[13] , \B_DOUT_TEMPR96[13] , 
        \B_DOUT_TEMPR97[13] , \B_DOUT_TEMPR98[13] , 
        \B_DOUT_TEMPR99[13] , \B_DOUT_TEMPR100[13] , 
        \B_DOUT_TEMPR101[13] , \B_DOUT_TEMPR102[13] , 
        \B_DOUT_TEMPR103[13] , \B_DOUT_TEMPR104[13] , 
        \B_DOUT_TEMPR105[13] , \B_DOUT_TEMPR106[13] , 
        \B_DOUT_TEMPR107[13] , \B_DOUT_TEMPR108[13] , 
        \B_DOUT_TEMPR109[13] , \B_DOUT_TEMPR110[13] , 
        \B_DOUT_TEMPR111[13] , \B_DOUT_TEMPR112[13] , 
        \B_DOUT_TEMPR113[13] , \B_DOUT_TEMPR114[13] , 
        \B_DOUT_TEMPR115[13] , \B_DOUT_TEMPR116[13] , 
        \B_DOUT_TEMPR117[13] , \B_DOUT_TEMPR118[13] , 
        \B_DOUT_TEMPR0[14] , \B_DOUT_TEMPR1[14] , \B_DOUT_TEMPR2[14] , 
        \B_DOUT_TEMPR3[14] , \B_DOUT_TEMPR4[14] , \B_DOUT_TEMPR5[14] , 
        \B_DOUT_TEMPR6[14] , \B_DOUT_TEMPR7[14] , \B_DOUT_TEMPR8[14] , 
        \B_DOUT_TEMPR9[14] , \B_DOUT_TEMPR10[14] , 
        \B_DOUT_TEMPR11[14] , \B_DOUT_TEMPR12[14] , 
        \B_DOUT_TEMPR13[14] , \B_DOUT_TEMPR14[14] , 
        \B_DOUT_TEMPR15[14] , \B_DOUT_TEMPR16[14] , 
        \B_DOUT_TEMPR17[14] , \B_DOUT_TEMPR18[14] , 
        \B_DOUT_TEMPR19[14] , \B_DOUT_TEMPR20[14] , 
        \B_DOUT_TEMPR21[14] , \B_DOUT_TEMPR22[14] , 
        \B_DOUT_TEMPR23[14] , \B_DOUT_TEMPR24[14] , 
        \B_DOUT_TEMPR25[14] , \B_DOUT_TEMPR26[14] , 
        \B_DOUT_TEMPR27[14] , \B_DOUT_TEMPR28[14] , 
        \B_DOUT_TEMPR29[14] , \B_DOUT_TEMPR30[14] , 
        \B_DOUT_TEMPR31[14] , \B_DOUT_TEMPR32[14] , 
        \B_DOUT_TEMPR33[14] , \B_DOUT_TEMPR34[14] , 
        \B_DOUT_TEMPR35[14] , \B_DOUT_TEMPR36[14] , 
        \B_DOUT_TEMPR37[14] , \B_DOUT_TEMPR38[14] , 
        \B_DOUT_TEMPR39[14] , \B_DOUT_TEMPR40[14] , 
        \B_DOUT_TEMPR41[14] , \B_DOUT_TEMPR42[14] , 
        \B_DOUT_TEMPR43[14] , \B_DOUT_TEMPR44[14] , 
        \B_DOUT_TEMPR45[14] , \B_DOUT_TEMPR46[14] , 
        \B_DOUT_TEMPR47[14] , \B_DOUT_TEMPR48[14] , 
        \B_DOUT_TEMPR49[14] , \B_DOUT_TEMPR50[14] , 
        \B_DOUT_TEMPR51[14] , \B_DOUT_TEMPR52[14] , 
        \B_DOUT_TEMPR53[14] , \B_DOUT_TEMPR54[14] , 
        \B_DOUT_TEMPR55[14] , \B_DOUT_TEMPR56[14] , 
        \B_DOUT_TEMPR57[14] , \B_DOUT_TEMPR58[14] , 
        \B_DOUT_TEMPR59[14] , \B_DOUT_TEMPR60[14] , 
        \B_DOUT_TEMPR61[14] , \B_DOUT_TEMPR62[14] , 
        \B_DOUT_TEMPR63[14] , \B_DOUT_TEMPR64[14] , 
        \B_DOUT_TEMPR65[14] , \B_DOUT_TEMPR66[14] , 
        \B_DOUT_TEMPR67[14] , \B_DOUT_TEMPR68[14] , 
        \B_DOUT_TEMPR69[14] , \B_DOUT_TEMPR70[14] , 
        \B_DOUT_TEMPR71[14] , \B_DOUT_TEMPR72[14] , 
        \B_DOUT_TEMPR73[14] , \B_DOUT_TEMPR74[14] , 
        \B_DOUT_TEMPR75[14] , \B_DOUT_TEMPR76[14] , 
        \B_DOUT_TEMPR77[14] , \B_DOUT_TEMPR78[14] , 
        \B_DOUT_TEMPR79[14] , \B_DOUT_TEMPR80[14] , 
        \B_DOUT_TEMPR81[14] , \B_DOUT_TEMPR82[14] , 
        \B_DOUT_TEMPR83[14] , \B_DOUT_TEMPR84[14] , 
        \B_DOUT_TEMPR85[14] , \B_DOUT_TEMPR86[14] , 
        \B_DOUT_TEMPR87[14] , \B_DOUT_TEMPR88[14] , 
        \B_DOUT_TEMPR89[14] , \B_DOUT_TEMPR90[14] , 
        \B_DOUT_TEMPR91[14] , \B_DOUT_TEMPR92[14] , 
        \B_DOUT_TEMPR93[14] , \B_DOUT_TEMPR94[14] , 
        \B_DOUT_TEMPR95[14] , \B_DOUT_TEMPR96[14] , 
        \B_DOUT_TEMPR97[14] , \B_DOUT_TEMPR98[14] , 
        \B_DOUT_TEMPR99[14] , \B_DOUT_TEMPR100[14] , 
        \B_DOUT_TEMPR101[14] , \B_DOUT_TEMPR102[14] , 
        \B_DOUT_TEMPR103[14] , \B_DOUT_TEMPR104[14] , 
        \B_DOUT_TEMPR105[14] , \B_DOUT_TEMPR106[14] , 
        \B_DOUT_TEMPR107[14] , \B_DOUT_TEMPR108[14] , 
        \B_DOUT_TEMPR109[14] , \B_DOUT_TEMPR110[14] , 
        \B_DOUT_TEMPR111[14] , \B_DOUT_TEMPR112[14] , 
        \B_DOUT_TEMPR113[14] , \B_DOUT_TEMPR114[14] , 
        \B_DOUT_TEMPR115[14] , \B_DOUT_TEMPR116[14] , 
        \B_DOUT_TEMPR117[14] , \B_DOUT_TEMPR118[14] , 
        \B_DOUT_TEMPR0[15] , \B_DOUT_TEMPR1[15] , \B_DOUT_TEMPR2[15] , 
        \B_DOUT_TEMPR3[15] , \B_DOUT_TEMPR4[15] , \B_DOUT_TEMPR5[15] , 
        \B_DOUT_TEMPR6[15] , \B_DOUT_TEMPR7[15] , \B_DOUT_TEMPR8[15] , 
        \B_DOUT_TEMPR9[15] , \B_DOUT_TEMPR10[15] , 
        \B_DOUT_TEMPR11[15] , \B_DOUT_TEMPR12[15] , 
        \B_DOUT_TEMPR13[15] , \B_DOUT_TEMPR14[15] , 
        \B_DOUT_TEMPR15[15] , \B_DOUT_TEMPR16[15] , 
        \B_DOUT_TEMPR17[15] , \B_DOUT_TEMPR18[15] , 
        \B_DOUT_TEMPR19[15] , \B_DOUT_TEMPR20[15] , 
        \B_DOUT_TEMPR21[15] , \B_DOUT_TEMPR22[15] , 
        \B_DOUT_TEMPR23[15] , \B_DOUT_TEMPR24[15] , 
        \B_DOUT_TEMPR25[15] , \B_DOUT_TEMPR26[15] , 
        \B_DOUT_TEMPR27[15] , \B_DOUT_TEMPR28[15] , 
        \B_DOUT_TEMPR29[15] , \B_DOUT_TEMPR30[15] , 
        \B_DOUT_TEMPR31[15] , \B_DOUT_TEMPR32[15] , 
        \B_DOUT_TEMPR33[15] , \B_DOUT_TEMPR34[15] , 
        \B_DOUT_TEMPR35[15] , \B_DOUT_TEMPR36[15] , 
        \B_DOUT_TEMPR37[15] , \B_DOUT_TEMPR38[15] , 
        \B_DOUT_TEMPR39[15] , \B_DOUT_TEMPR40[15] , 
        \B_DOUT_TEMPR41[15] , \B_DOUT_TEMPR42[15] , 
        \B_DOUT_TEMPR43[15] , \B_DOUT_TEMPR44[15] , 
        \B_DOUT_TEMPR45[15] , \B_DOUT_TEMPR46[15] , 
        \B_DOUT_TEMPR47[15] , \B_DOUT_TEMPR48[15] , 
        \B_DOUT_TEMPR49[15] , \B_DOUT_TEMPR50[15] , 
        \B_DOUT_TEMPR51[15] , \B_DOUT_TEMPR52[15] , 
        \B_DOUT_TEMPR53[15] , \B_DOUT_TEMPR54[15] , 
        \B_DOUT_TEMPR55[15] , \B_DOUT_TEMPR56[15] , 
        \B_DOUT_TEMPR57[15] , \B_DOUT_TEMPR58[15] , 
        \B_DOUT_TEMPR59[15] , \B_DOUT_TEMPR60[15] , 
        \B_DOUT_TEMPR61[15] , \B_DOUT_TEMPR62[15] , 
        \B_DOUT_TEMPR63[15] , \B_DOUT_TEMPR64[15] , 
        \B_DOUT_TEMPR65[15] , \B_DOUT_TEMPR66[15] , 
        \B_DOUT_TEMPR67[15] , \B_DOUT_TEMPR68[15] , 
        \B_DOUT_TEMPR69[15] , \B_DOUT_TEMPR70[15] , 
        \B_DOUT_TEMPR71[15] , \B_DOUT_TEMPR72[15] , 
        \B_DOUT_TEMPR73[15] , \B_DOUT_TEMPR74[15] , 
        \B_DOUT_TEMPR75[15] , \B_DOUT_TEMPR76[15] , 
        \B_DOUT_TEMPR77[15] , \B_DOUT_TEMPR78[15] , 
        \B_DOUT_TEMPR79[15] , \B_DOUT_TEMPR80[15] , 
        \B_DOUT_TEMPR81[15] , \B_DOUT_TEMPR82[15] , 
        \B_DOUT_TEMPR83[15] , \B_DOUT_TEMPR84[15] , 
        \B_DOUT_TEMPR85[15] , \B_DOUT_TEMPR86[15] , 
        \B_DOUT_TEMPR87[15] , \B_DOUT_TEMPR88[15] , 
        \B_DOUT_TEMPR89[15] , \B_DOUT_TEMPR90[15] , 
        \B_DOUT_TEMPR91[15] , \B_DOUT_TEMPR92[15] , 
        \B_DOUT_TEMPR93[15] , \B_DOUT_TEMPR94[15] , 
        \B_DOUT_TEMPR95[15] , \B_DOUT_TEMPR96[15] , 
        \B_DOUT_TEMPR97[15] , \B_DOUT_TEMPR98[15] , 
        \B_DOUT_TEMPR99[15] , \B_DOUT_TEMPR100[15] , 
        \B_DOUT_TEMPR101[15] , \B_DOUT_TEMPR102[15] , 
        \B_DOUT_TEMPR103[15] , \B_DOUT_TEMPR104[15] , 
        \B_DOUT_TEMPR105[15] , \B_DOUT_TEMPR106[15] , 
        \B_DOUT_TEMPR107[15] , \B_DOUT_TEMPR108[15] , 
        \B_DOUT_TEMPR109[15] , \B_DOUT_TEMPR110[15] , 
        \B_DOUT_TEMPR111[15] , \B_DOUT_TEMPR112[15] , 
        \B_DOUT_TEMPR113[15] , \B_DOUT_TEMPR114[15] , 
        \B_DOUT_TEMPR115[15] , \B_DOUT_TEMPR116[15] , 
        \B_DOUT_TEMPR117[15] , \B_DOUT_TEMPR118[15] , 
        \B_DOUT_TEMPR0[16] , \B_DOUT_TEMPR1[16] , \B_DOUT_TEMPR2[16] , 
        \B_DOUT_TEMPR3[16] , \B_DOUT_TEMPR4[16] , \B_DOUT_TEMPR5[16] , 
        \B_DOUT_TEMPR6[16] , \B_DOUT_TEMPR7[16] , \B_DOUT_TEMPR8[16] , 
        \B_DOUT_TEMPR9[16] , \B_DOUT_TEMPR10[16] , 
        \B_DOUT_TEMPR11[16] , \B_DOUT_TEMPR12[16] , 
        \B_DOUT_TEMPR13[16] , \B_DOUT_TEMPR14[16] , 
        \B_DOUT_TEMPR15[16] , \B_DOUT_TEMPR16[16] , 
        \B_DOUT_TEMPR17[16] , \B_DOUT_TEMPR18[16] , 
        \B_DOUT_TEMPR19[16] , \B_DOUT_TEMPR20[16] , 
        \B_DOUT_TEMPR21[16] , \B_DOUT_TEMPR22[16] , 
        \B_DOUT_TEMPR23[16] , \B_DOUT_TEMPR24[16] , 
        \B_DOUT_TEMPR25[16] , \B_DOUT_TEMPR26[16] , 
        \B_DOUT_TEMPR27[16] , \B_DOUT_TEMPR28[16] , 
        \B_DOUT_TEMPR29[16] , \B_DOUT_TEMPR30[16] , 
        \B_DOUT_TEMPR31[16] , \B_DOUT_TEMPR32[16] , 
        \B_DOUT_TEMPR33[16] , \B_DOUT_TEMPR34[16] , 
        \B_DOUT_TEMPR35[16] , \B_DOUT_TEMPR36[16] , 
        \B_DOUT_TEMPR37[16] , \B_DOUT_TEMPR38[16] , 
        \B_DOUT_TEMPR39[16] , \B_DOUT_TEMPR40[16] , 
        \B_DOUT_TEMPR41[16] , \B_DOUT_TEMPR42[16] , 
        \B_DOUT_TEMPR43[16] , \B_DOUT_TEMPR44[16] , 
        \B_DOUT_TEMPR45[16] , \B_DOUT_TEMPR46[16] , 
        \B_DOUT_TEMPR47[16] , \B_DOUT_TEMPR48[16] , 
        \B_DOUT_TEMPR49[16] , \B_DOUT_TEMPR50[16] , 
        \B_DOUT_TEMPR51[16] , \B_DOUT_TEMPR52[16] , 
        \B_DOUT_TEMPR53[16] , \B_DOUT_TEMPR54[16] , 
        \B_DOUT_TEMPR55[16] , \B_DOUT_TEMPR56[16] , 
        \B_DOUT_TEMPR57[16] , \B_DOUT_TEMPR58[16] , 
        \B_DOUT_TEMPR59[16] , \B_DOUT_TEMPR60[16] , 
        \B_DOUT_TEMPR61[16] , \B_DOUT_TEMPR62[16] , 
        \B_DOUT_TEMPR63[16] , \B_DOUT_TEMPR64[16] , 
        \B_DOUT_TEMPR65[16] , \B_DOUT_TEMPR66[16] , 
        \B_DOUT_TEMPR67[16] , \B_DOUT_TEMPR68[16] , 
        \B_DOUT_TEMPR69[16] , \B_DOUT_TEMPR70[16] , 
        \B_DOUT_TEMPR71[16] , \B_DOUT_TEMPR72[16] , 
        \B_DOUT_TEMPR73[16] , \B_DOUT_TEMPR74[16] , 
        \B_DOUT_TEMPR75[16] , \B_DOUT_TEMPR76[16] , 
        \B_DOUT_TEMPR77[16] , \B_DOUT_TEMPR78[16] , 
        \B_DOUT_TEMPR79[16] , \B_DOUT_TEMPR80[16] , 
        \B_DOUT_TEMPR81[16] , \B_DOUT_TEMPR82[16] , 
        \B_DOUT_TEMPR83[16] , \B_DOUT_TEMPR84[16] , 
        \B_DOUT_TEMPR85[16] , \B_DOUT_TEMPR86[16] , 
        \B_DOUT_TEMPR87[16] , \B_DOUT_TEMPR88[16] , 
        \B_DOUT_TEMPR89[16] , \B_DOUT_TEMPR90[16] , 
        \B_DOUT_TEMPR91[16] , \B_DOUT_TEMPR92[16] , 
        \B_DOUT_TEMPR93[16] , \B_DOUT_TEMPR94[16] , 
        \B_DOUT_TEMPR95[16] , \B_DOUT_TEMPR96[16] , 
        \B_DOUT_TEMPR97[16] , \B_DOUT_TEMPR98[16] , 
        \B_DOUT_TEMPR99[16] , \B_DOUT_TEMPR100[16] , 
        \B_DOUT_TEMPR101[16] , \B_DOUT_TEMPR102[16] , 
        \B_DOUT_TEMPR103[16] , \B_DOUT_TEMPR104[16] , 
        \B_DOUT_TEMPR105[16] , \B_DOUT_TEMPR106[16] , 
        \B_DOUT_TEMPR107[16] , \B_DOUT_TEMPR108[16] , 
        \B_DOUT_TEMPR109[16] , \B_DOUT_TEMPR110[16] , 
        \B_DOUT_TEMPR111[16] , \B_DOUT_TEMPR112[16] , 
        \B_DOUT_TEMPR113[16] , \B_DOUT_TEMPR114[16] , 
        \B_DOUT_TEMPR115[16] , \B_DOUT_TEMPR116[16] , 
        \B_DOUT_TEMPR117[16] , \B_DOUT_TEMPR118[16] , 
        \B_DOUT_TEMPR0[17] , \B_DOUT_TEMPR1[17] , \B_DOUT_TEMPR2[17] , 
        \B_DOUT_TEMPR3[17] , \B_DOUT_TEMPR4[17] , \B_DOUT_TEMPR5[17] , 
        \B_DOUT_TEMPR6[17] , \B_DOUT_TEMPR7[17] , \B_DOUT_TEMPR8[17] , 
        \B_DOUT_TEMPR9[17] , \B_DOUT_TEMPR10[17] , 
        \B_DOUT_TEMPR11[17] , \B_DOUT_TEMPR12[17] , 
        \B_DOUT_TEMPR13[17] , \B_DOUT_TEMPR14[17] , 
        \B_DOUT_TEMPR15[17] , \B_DOUT_TEMPR16[17] , 
        \B_DOUT_TEMPR17[17] , \B_DOUT_TEMPR18[17] , 
        \B_DOUT_TEMPR19[17] , \B_DOUT_TEMPR20[17] , 
        \B_DOUT_TEMPR21[17] , \B_DOUT_TEMPR22[17] , 
        \B_DOUT_TEMPR23[17] , \B_DOUT_TEMPR24[17] , 
        \B_DOUT_TEMPR25[17] , \B_DOUT_TEMPR26[17] , 
        \B_DOUT_TEMPR27[17] , \B_DOUT_TEMPR28[17] , 
        \B_DOUT_TEMPR29[17] , \B_DOUT_TEMPR30[17] , 
        \B_DOUT_TEMPR31[17] , \B_DOUT_TEMPR32[17] , 
        \B_DOUT_TEMPR33[17] , \B_DOUT_TEMPR34[17] , 
        \B_DOUT_TEMPR35[17] , \B_DOUT_TEMPR36[17] , 
        \B_DOUT_TEMPR37[17] , \B_DOUT_TEMPR38[17] , 
        \B_DOUT_TEMPR39[17] , \B_DOUT_TEMPR40[17] , 
        \B_DOUT_TEMPR41[17] , \B_DOUT_TEMPR42[17] , 
        \B_DOUT_TEMPR43[17] , \B_DOUT_TEMPR44[17] , 
        \B_DOUT_TEMPR45[17] , \B_DOUT_TEMPR46[17] , 
        \B_DOUT_TEMPR47[17] , \B_DOUT_TEMPR48[17] , 
        \B_DOUT_TEMPR49[17] , \B_DOUT_TEMPR50[17] , 
        \B_DOUT_TEMPR51[17] , \B_DOUT_TEMPR52[17] , 
        \B_DOUT_TEMPR53[17] , \B_DOUT_TEMPR54[17] , 
        \B_DOUT_TEMPR55[17] , \B_DOUT_TEMPR56[17] , 
        \B_DOUT_TEMPR57[17] , \B_DOUT_TEMPR58[17] , 
        \B_DOUT_TEMPR59[17] , \B_DOUT_TEMPR60[17] , 
        \B_DOUT_TEMPR61[17] , \B_DOUT_TEMPR62[17] , 
        \B_DOUT_TEMPR63[17] , \B_DOUT_TEMPR64[17] , 
        \B_DOUT_TEMPR65[17] , \B_DOUT_TEMPR66[17] , 
        \B_DOUT_TEMPR67[17] , \B_DOUT_TEMPR68[17] , 
        \B_DOUT_TEMPR69[17] , \B_DOUT_TEMPR70[17] , 
        \B_DOUT_TEMPR71[17] , \B_DOUT_TEMPR72[17] , 
        \B_DOUT_TEMPR73[17] , \B_DOUT_TEMPR74[17] , 
        \B_DOUT_TEMPR75[17] , \B_DOUT_TEMPR76[17] , 
        \B_DOUT_TEMPR77[17] , \B_DOUT_TEMPR78[17] , 
        \B_DOUT_TEMPR79[17] , \B_DOUT_TEMPR80[17] , 
        \B_DOUT_TEMPR81[17] , \B_DOUT_TEMPR82[17] , 
        \B_DOUT_TEMPR83[17] , \B_DOUT_TEMPR84[17] , 
        \B_DOUT_TEMPR85[17] , \B_DOUT_TEMPR86[17] , 
        \B_DOUT_TEMPR87[17] , \B_DOUT_TEMPR88[17] , 
        \B_DOUT_TEMPR89[17] , \B_DOUT_TEMPR90[17] , 
        \B_DOUT_TEMPR91[17] , \B_DOUT_TEMPR92[17] , 
        \B_DOUT_TEMPR93[17] , \B_DOUT_TEMPR94[17] , 
        \B_DOUT_TEMPR95[17] , \B_DOUT_TEMPR96[17] , 
        \B_DOUT_TEMPR97[17] , \B_DOUT_TEMPR98[17] , 
        \B_DOUT_TEMPR99[17] , \B_DOUT_TEMPR100[17] , 
        \B_DOUT_TEMPR101[17] , \B_DOUT_TEMPR102[17] , 
        \B_DOUT_TEMPR103[17] , \B_DOUT_TEMPR104[17] , 
        \B_DOUT_TEMPR105[17] , \B_DOUT_TEMPR106[17] , 
        \B_DOUT_TEMPR107[17] , \B_DOUT_TEMPR108[17] , 
        \B_DOUT_TEMPR109[17] , \B_DOUT_TEMPR110[17] , 
        \B_DOUT_TEMPR111[17] , \B_DOUT_TEMPR112[17] , 
        \B_DOUT_TEMPR113[17] , \B_DOUT_TEMPR114[17] , 
        \B_DOUT_TEMPR115[17] , \B_DOUT_TEMPR116[17] , 
        \B_DOUT_TEMPR117[17] , \B_DOUT_TEMPR118[17] , 
        \B_DOUT_TEMPR0[18] , \B_DOUT_TEMPR1[18] , \B_DOUT_TEMPR2[18] , 
        \B_DOUT_TEMPR3[18] , \B_DOUT_TEMPR4[18] , \B_DOUT_TEMPR5[18] , 
        \B_DOUT_TEMPR6[18] , \B_DOUT_TEMPR7[18] , \B_DOUT_TEMPR8[18] , 
        \B_DOUT_TEMPR9[18] , \B_DOUT_TEMPR10[18] , 
        \B_DOUT_TEMPR11[18] , \B_DOUT_TEMPR12[18] , 
        \B_DOUT_TEMPR13[18] , \B_DOUT_TEMPR14[18] , 
        \B_DOUT_TEMPR15[18] , \B_DOUT_TEMPR16[18] , 
        \B_DOUT_TEMPR17[18] , \B_DOUT_TEMPR18[18] , 
        \B_DOUT_TEMPR19[18] , \B_DOUT_TEMPR20[18] , 
        \B_DOUT_TEMPR21[18] , \B_DOUT_TEMPR22[18] , 
        \B_DOUT_TEMPR23[18] , \B_DOUT_TEMPR24[18] , 
        \B_DOUT_TEMPR25[18] , \B_DOUT_TEMPR26[18] , 
        \B_DOUT_TEMPR27[18] , \B_DOUT_TEMPR28[18] , 
        \B_DOUT_TEMPR29[18] , \B_DOUT_TEMPR30[18] , 
        \B_DOUT_TEMPR31[18] , \B_DOUT_TEMPR32[18] , 
        \B_DOUT_TEMPR33[18] , \B_DOUT_TEMPR34[18] , 
        \B_DOUT_TEMPR35[18] , \B_DOUT_TEMPR36[18] , 
        \B_DOUT_TEMPR37[18] , \B_DOUT_TEMPR38[18] , 
        \B_DOUT_TEMPR39[18] , \B_DOUT_TEMPR40[18] , 
        \B_DOUT_TEMPR41[18] , \B_DOUT_TEMPR42[18] , 
        \B_DOUT_TEMPR43[18] , \B_DOUT_TEMPR44[18] , 
        \B_DOUT_TEMPR45[18] , \B_DOUT_TEMPR46[18] , 
        \B_DOUT_TEMPR47[18] , \B_DOUT_TEMPR48[18] , 
        \B_DOUT_TEMPR49[18] , \B_DOUT_TEMPR50[18] , 
        \B_DOUT_TEMPR51[18] , \B_DOUT_TEMPR52[18] , 
        \B_DOUT_TEMPR53[18] , \B_DOUT_TEMPR54[18] , 
        \B_DOUT_TEMPR55[18] , \B_DOUT_TEMPR56[18] , 
        \B_DOUT_TEMPR57[18] , \B_DOUT_TEMPR58[18] , 
        \B_DOUT_TEMPR59[18] , \B_DOUT_TEMPR60[18] , 
        \B_DOUT_TEMPR61[18] , \B_DOUT_TEMPR62[18] , 
        \B_DOUT_TEMPR63[18] , \B_DOUT_TEMPR64[18] , 
        \B_DOUT_TEMPR65[18] , \B_DOUT_TEMPR66[18] , 
        \B_DOUT_TEMPR67[18] , \B_DOUT_TEMPR68[18] , 
        \B_DOUT_TEMPR69[18] , \B_DOUT_TEMPR70[18] , 
        \B_DOUT_TEMPR71[18] , \B_DOUT_TEMPR72[18] , 
        \B_DOUT_TEMPR73[18] , \B_DOUT_TEMPR74[18] , 
        \B_DOUT_TEMPR75[18] , \B_DOUT_TEMPR76[18] , 
        \B_DOUT_TEMPR77[18] , \B_DOUT_TEMPR78[18] , 
        \B_DOUT_TEMPR79[18] , \B_DOUT_TEMPR80[18] , 
        \B_DOUT_TEMPR81[18] , \B_DOUT_TEMPR82[18] , 
        \B_DOUT_TEMPR83[18] , \B_DOUT_TEMPR84[18] , 
        \B_DOUT_TEMPR85[18] , \B_DOUT_TEMPR86[18] , 
        \B_DOUT_TEMPR87[18] , \B_DOUT_TEMPR88[18] , 
        \B_DOUT_TEMPR89[18] , \B_DOUT_TEMPR90[18] , 
        \B_DOUT_TEMPR91[18] , \B_DOUT_TEMPR92[18] , 
        \B_DOUT_TEMPR93[18] , \B_DOUT_TEMPR94[18] , 
        \B_DOUT_TEMPR95[18] , \B_DOUT_TEMPR96[18] , 
        \B_DOUT_TEMPR97[18] , \B_DOUT_TEMPR98[18] , 
        \B_DOUT_TEMPR99[18] , \B_DOUT_TEMPR100[18] , 
        \B_DOUT_TEMPR101[18] , \B_DOUT_TEMPR102[18] , 
        \B_DOUT_TEMPR103[18] , \B_DOUT_TEMPR104[18] , 
        \B_DOUT_TEMPR105[18] , \B_DOUT_TEMPR106[18] , 
        \B_DOUT_TEMPR107[18] , \B_DOUT_TEMPR108[18] , 
        \B_DOUT_TEMPR109[18] , \B_DOUT_TEMPR110[18] , 
        \B_DOUT_TEMPR111[18] , \B_DOUT_TEMPR112[18] , 
        \B_DOUT_TEMPR113[18] , \B_DOUT_TEMPR114[18] , 
        \B_DOUT_TEMPR115[18] , \B_DOUT_TEMPR116[18] , 
        \B_DOUT_TEMPR117[18] , \B_DOUT_TEMPR118[18] , 
        \B_DOUT_TEMPR0[19] , \B_DOUT_TEMPR1[19] , \B_DOUT_TEMPR2[19] , 
        \B_DOUT_TEMPR3[19] , \B_DOUT_TEMPR4[19] , \B_DOUT_TEMPR5[19] , 
        \B_DOUT_TEMPR6[19] , \B_DOUT_TEMPR7[19] , \B_DOUT_TEMPR8[19] , 
        \B_DOUT_TEMPR9[19] , \B_DOUT_TEMPR10[19] , 
        \B_DOUT_TEMPR11[19] , \B_DOUT_TEMPR12[19] , 
        \B_DOUT_TEMPR13[19] , \B_DOUT_TEMPR14[19] , 
        \B_DOUT_TEMPR15[19] , \B_DOUT_TEMPR16[19] , 
        \B_DOUT_TEMPR17[19] , \B_DOUT_TEMPR18[19] , 
        \B_DOUT_TEMPR19[19] , \B_DOUT_TEMPR20[19] , 
        \B_DOUT_TEMPR21[19] , \B_DOUT_TEMPR22[19] , 
        \B_DOUT_TEMPR23[19] , \B_DOUT_TEMPR24[19] , 
        \B_DOUT_TEMPR25[19] , \B_DOUT_TEMPR26[19] , 
        \B_DOUT_TEMPR27[19] , \B_DOUT_TEMPR28[19] , 
        \B_DOUT_TEMPR29[19] , \B_DOUT_TEMPR30[19] , 
        \B_DOUT_TEMPR31[19] , \B_DOUT_TEMPR32[19] , 
        \B_DOUT_TEMPR33[19] , \B_DOUT_TEMPR34[19] , 
        \B_DOUT_TEMPR35[19] , \B_DOUT_TEMPR36[19] , 
        \B_DOUT_TEMPR37[19] , \B_DOUT_TEMPR38[19] , 
        \B_DOUT_TEMPR39[19] , \B_DOUT_TEMPR40[19] , 
        \B_DOUT_TEMPR41[19] , \B_DOUT_TEMPR42[19] , 
        \B_DOUT_TEMPR43[19] , \B_DOUT_TEMPR44[19] , 
        \B_DOUT_TEMPR45[19] , \B_DOUT_TEMPR46[19] , 
        \B_DOUT_TEMPR47[19] , \B_DOUT_TEMPR48[19] , 
        \B_DOUT_TEMPR49[19] , \B_DOUT_TEMPR50[19] , 
        \B_DOUT_TEMPR51[19] , \B_DOUT_TEMPR52[19] , 
        \B_DOUT_TEMPR53[19] , \B_DOUT_TEMPR54[19] , 
        \B_DOUT_TEMPR55[19] , \B_DOUT_TEMPR56[19] , 
        \B_DOUT_TEMPR57[19] , \B_DOUT_TEMPR58[19] , 
        \B_DOUT_TEMPR59[19] , \B_DOUT_TEMPR60[19] , 
        \B_DOUT_TEMPR61[19] , \B_DOUT_TEMPR62[19] , 
        \B_DOUT_TEMPR63[19] , \B_DOUT_TEMPR64[19] , 
        \B_DOUT_TEMPR65[19] , \B_DOUT_TEMPR66[19] , 
        \B_DOUT_TEMPR67[19] , \B_DOUT_TEMPR68[19] , 
        \B_DOUT_TEMPR69[19] , \B_DOUT_TEMPR70[19] , 
        \B_DOUT_TEMPR71[19] , \B_DOUT_TEMPR72[19] , 
        \B_DOUT_TEMPR73[19] , \B_DOUT_TEMPR74[19] , 
        \B_DOUT_TEMPR75[19] , \B_DOUT_TEMPR76[19] , 
        \B_DOUT_TEMPR77[19] , \B_DOUT_TEMPR78[19] , 
        \B_DOUT_TEMPR79[19] , \B_DOUT_TEMPR80[19] , 
        \B_DOUT_TEMPR81[19] , \B_DOUT_TEMPR82[19] , 
        \B_DOUT_TEMPR83[19] , \B_DOUT_TEMPR84[19] , 
        \B_DOUT_TEMPR85[19] , \B_DOUT_TEMPR86[19] , 
        \B_DOUT_TEMPR87[19] , \B_DOUT_TEMPR88[19] , 
        \B_DOUT_TEMPR89[19] , \B_DOUT_TEMPR90[19] , 
        \B_DOUT_TEMPR91[19] , \B_DOUT_TEMPR92[19] , 
        \B_DOUT_TEMPR93[19] , \B_DOUT_TEMPR94[19] , 
        \B_DOUT_TEMPR95[19] , \B_DOUT_TEMPR96[19] , 
        \B_DOUT_TEMPR97[19] , \B_DOUT_TEMPR98[19] , 
        \B_DOUT_TEMPR99[19] , \B_DOUT_TEMPR100[19] , 
        \B_DOUT_TEMPR101[19] , \B_DOUT_TEMPR102[19] , 
        \B_DOUT_TEMPR103[19] , \B_DOUT_TEMPR104[19] , 
        \B_DOUT_TEMPR105[19] , \B_DOUT_TEMPR106[19] , 
        \B_DOUT_TEMPR107[19] , \B_DOUT_TEMPR108[19] , 
        \B_DOUT_TEMPR109[19] , \B_DOUT_TEMPR110[19] , 
        \B_DOUT_TEMPR111[19] , \B_DOUT_TEMPR112[19] , 
        \B_DOUT_TEMPR113[19] , \B_DOUT_TEMPR114[19] , 
        \B_DOUT_TEMPR115[19] , \B_DOUT_TEMPR116[19] , 
        \B_DOUT_TEMPR117[19] , \B_DOUT_TEMPR118[19] , 
        \B_DOUT_TEMPR0[20] , \B_DOUT_TEMPR1[20] , \B_DOUT_TEMPR2[20] , 
        \B_DOUT_TEMPR3[20] , \B_DOUT_TEMPR4[20] , \B_DOUT_TEMPR5[20] , 
        \B_DOUT_TEMPR6[20] , \B_DOUT_TEMPR7[20] , \B_DOUT_TEMPR8[20] , 
        \B_DOUT_TEMPR9[20] , \B_DOUT_TEMPR10[20] , 
        \B_DOUT_TEMPR11[20] , \B_DOUT_TEMPR12[20] , 
        \B_DOUT_TEMPR13[20] , \B_DOUT_TEMPR14[20] , 
        \B_DOUT_TEMPR15[20] , \B_DOUT_TEMPR16[20] , 
        \B_DOUT_TEMPR17[20] , \B_DOUT_TEMPR18[20] , 
        \B_DOUT_TEMPR19[20] , \B_DOUT_TEMPR20[20] , 
        \B_DOUT_TEMPR21[20] , \B_DOUT_TEMPR22[20] , 
        \B_DOUT_TEMPR23[20] , \B_DOUT_TEMPR24[20] , 
        \B_DOUT_TEMPR25[20] , \B_DOUT_TEMPR26[20] , 
        \B_DOUT_TEMPR27[20] , \B_DOUT_TEMPR28[20] , 
        \B_DOUT_TEMPR29[20] , \B_DOUT_TEMPR30[20] , 
        \B_DOUT_TEMPR31[20] , \B_DOUT_TEMPR32[20] , 
        \B_DOUT_TEMPR33[20] , \B_DOUT_TEMPR34[20] , 
        \B_DOUT_TEMPR35[20] , \B_DOUT_TEMPR36[20] , 
        \B_DOUT_TEMPR37[20] , \B_DOUT_TEMPR38[20] , 
        \B_DOUT_TEMPR39[20] , \B_DOUT_TEMPR40[20] , 
        \B_DOUT_TEMPR41[20] , \B_DOUT_TEMPR42[20] , 
        \B_DOUT_TEMPR43[20] , \B_DOUT_TEMPR44[20] , 
        \B_DOUT_TEMPR45[20] , \B_DOUT_TEMPR46[20] , 
        \B_DOUT_TEMPR47[20] , \B_DOUT_TEMPR48[20] , 
        \B_DOUT_TEMPR49[20] , \B_DOUT_TEMPR50[20] , 
        \B_DOUT_TEMPR51[20] , \B_DOUT_TEMPR52[20] , 
        \B_DOUT_TEMPR53[20] , \B_DOUT_TEMPR54[20] , 
        \B_DOUT_TEMPR55[20] , \B_DOUT_TEMPR56[20] , 
        \B_DOUT_TEMPR57[20] , \B_DOUT_TEMPR58[20] , 
        \B_DOUT_TEMPR59[20] , \B_DOUT_TEMPR60[20] , 
        \B_DOUT_TEMPR61[20] , \B_DOUT_TEMPR62[20] , 
        \B_DOUT_TEMPR63[20] , \B_DOUT_TEMPR64[20] , 
        \B_DOUT_TEMPR65[20] , \B_DOUT_TEMPR66[20] , 
        \B_DOUT_TEMPR67[20] , \B_DOUT_TEMPR68[20] , 
        \B_DOUT_TEMPR69[20] , \B_DOUT_TEMPR70[20] , 
        \B_DOUT_TEMPR71[20] , \B_DOUT_TEMPR72[20] , 
        \B_DOUT_TEMPR73[20] , \B_DOUT_TEMPR74[20] , 
        \B_DOUT_TEMPR75[20] , \B_DOUT_TEMPR76[20] , 
        \B_DOUT_TEMPR77[20] , \B_DOUT_TEMPR78[20] , 
        \B_DOUT_TEMPR79[20] , \B_DOUT_TEMPR80[20] , 
        \B_DOUT_TEMPR81[20] , \B_DOUT_TEMPR82[20] , 
        \B_DOUT_TEMPR83[20] , \B_DOUT_TEMPR84[20] , 
        \B_DOUT_TEMPR85[20] , \B_DOUT_TEMPR86[20] , 
        \B_DOUT_TEMPR87[20] , \B_DOUT_TEMPR88[20] , 
        \B_DOUT_TEMPR89[20] , \B_DOUT_TEMPR90[20] , 
        \B_DOUT_TEMPR91[20] , \B_DOUT_TEMPR92[20] , 
        \B_DOUT_TEMPR93[20] , \B_DOUT_TEMPR94[20] , 
        \B_DOUT_TEMPR95[20] , \B_DOUT_TEMPR96[20] , 
        \B_DOUT_TEMPR97[20] , \B_DOUT_TEMPR98[20] , 
        \B_DOUT_TEMPR99[20] , \B_DOUT_TEMPR100[20] , 
        \B_DOUT_TEMPR101[20] , \B_DOUT_TEMPR102[20] , 
        \B_DOUT_TEMPR103[20] , \B_DOUT_TEMPR104[20] , 
        \B_DOUT_TEMPR105[20] , \B_DOUT_TEMPR106[20] , 
        \B_DOUT_TEMPR107[20] , \B_DOUT_TEMPR108[20] , 
        \B_DOUT_TEMPR109[20] , \B_DOUT_TEMPR110[20] , 
        \B_DOUT_TEMPR111[20] , \B_DOUT_TEMPR112[20] , 
        \B_DOUT_TEMPR113[20] , \B_DOUT_TEMPR114[20] , 
        \B_DOUT_TEMPR115[20] , \B_DOUT_TEMPR116[20] , 
        \B_DOUT_TEMPR117[20] , \B_DOUT_TEMPR118[20] , 
        \B_DOUT_TEMPR0[21] , \B_DOUT_TEMPR1[21] , \B_DOUT_TEMPR2[21] , 
        \B_DOUT_TEMPR3[21] , \B_DOUT_TEMPR4[21] , \B_DOUT_TEMPR5[21] , 
        \B_DOUT_TEMPR6[21] , \B_DOUT_TEMPR7[21] , \B_DOUT_TEMPR8[21] , 
        \B_DOUT_TEMPR9[21] , \B_DOUT_TEMPR10[21] , 
        \B_DOUT_TEMPR11[21] , \B_DOUT_TEMPR12[21] , 
        \B_DOUT_TEMPR13[21] , \B_DOUT_TEMPR14[21] , 
        \B_DOUT_TEMPR15[21] , \B_DOUT_TEMPR16[21] , 
        \B_DOUT_TEMPR17[21] , \B_DOUT_TEMPR18[21] , 
        \B_DOUT_TEMPR19[21] , \B_DOUT_TEMPR20[21] , 
        \B_DOUT_TEMPR21[21] , \B_DOUT_TEMPR22[21] , 
        \B_DOUT_TEMPR23[21] , \B_DOUT_TEMPR24[21] , 
        \B_DOUT_TEMPR25[21] , \B_DOUT_TEMPR26[21] , 
        \B_DOUT_TEMPR27[21] , \B_DOUT_TEMPR28[21] , 
        \B_DOUT_TEMPR29[21] , \B_DOUT_TEMPR30[21] , 
        \B_DOUT_TEMPR31[21] , \B_DOUT_TEMPR32[21] , 
        \B_DOUT_TEMPR33[21] , \B_DOUT_TEMPR34[21] , 
        \B_DOUT_TEMPR35[21] , \B_DOUT_TEMPR36[21] , 
        \B_DOUT_TEMPR37[21] , \B_DOUT_TEMPR38[21] , 
        \B_DOUT_TEMPR39[21] , \B_DOUT_TEMPR40[21] , 
        \B_DOUT_TEMPR41[21] , \B_DOUT_TEMPR42[21] , 
        \B_DOUT_TEMPR43[21] , \B_DOUT_TEMPR44[21] , 
        \B_DOUT_TEMPR45[21] , \B_DOUT_TEMPR46[21] , 
        \B_DOUT_TEMPR47[21] , \B_DOUT_TEMPR48[21] , 
        \B_DOUT_TEMPR49[21] , \B_DOUT_TEMPR50[21] , 
        \B_DOUT_TEMPR51[21] , \B_DOUT_TEMPR52[21] , 
        \B_DOUT_TEMPR53[21] , \B_DOUT_TEMPR54[21] , 
        \B_DOUT_TEMPR55[21] , \B_DOUT_TEMPR56[21] , 
        \B_DOUT_TEMPR57[21] , \B_DOUT_TEMPR58[21] , 
        \B_DOUT_TEMPR59[21] , \B_DOUT_TEMPR60[21] , 
        \B_DOUT_TEMPR61[21] , \B_DOUT_TEMPR62[21] , 
        \B_DOUT_TEMPR63[21] , \B_DOUT_TEMPR64[21] , 
        \B_DOUT_TEMPR65[21] , \B_DOUT_TEMPR66[21] , 
        \B_DOUT_TEMPR67[21] , \B_DOUT_TEMPR68[21] , 
        \B_DOUT_TEMPR69[21] , \B_DOUT_TEMPR70[21] , 
        \B_DOUT_TEMPR71[21] , \B_DOUT_TEMPR72[21] , 
        \B_DOUT_TEMPR73[21] , \B_DOUT_TEMPR74[21] , 
        \B_DOUT_TEMPR75[21] , \B_DOUT_TEMPR76[21] , 
        \B_DOUT_TEMPR77[21] , \B_DOUT_TEMPR78[21] , 
        \B_DOUT_TEMPR79[21] , \B_DOUT_TEMPR80[21] , 
        \B_DOUT_TEMPR81[21] , \B_DOUT_TEMPR82[21] , 
        \B_DOUT_TEMPR83[21] , \B_DOUT_TEMPR84[21] , 
        \B_DOUT_TEMPR85[21] , \B_DOUT_TEMPR86[21] , 
        \B_DOUT_TEMPR87[21] , \B_DOUT_TEMPR88[21] , 
        \B_DOUT_TEMPR89[21] , \B_DOUT_TEMPR90[21] , 
        \B_DOUT_TEMPR91[21] , \B_DOUT_TEMPR92[21] , 
        \B_DOUT_TEMPR93[21] , \B_DOUT_TEMPR94[21] , 
        \B_DOUT_TEMPR95[21] , \B_DOUT_TEMPR96[21] , 
        \B_DOUT_TEMPR97[21] , \B_DOUT_TEMPR98[21] , 
        \B_DOUT_TEMPR99[21] , \B_DOUT_TEMPR100[21] , 
        \B_DOUT_TEMPR101[21] , \B_DOUT_TEMPR102[21] , 
        \B_DOUT_TEMPR103[21] , \B_DOUT_TEMPR104[21] , 
        \B_DOUT_TEMPR105[21] , \B_DOUT_TEMPR106[21] , 
        \B_DOUT_TEMPR107[21] , \B_DOUT_TEMPR108[21] , 
        \B_DOUT_TEMPR109[21] , \B_DOUT_TEMPR110[21] , 
        \B_DOUT_TEMPR111[21] , \B_DOUT_TEMPR112[21] , 
        \B_DOUT_TEMPR113[21] , \B_DOUT_TEMPR114[21] , 
        \B_DOUT_TEMPR115[21] , \B_DOUT_TEMPR116[21] , 
        \B_DOUT_TEMPR117[21] , \B_DOUT_TEMPR118[21] , 
        \B_DOUT_TEMPR0[22] , \B_DOUT_TEMPR1[22] , \B_DOUT_TEMPR2[22] , 
        \B_DOUT_TEMPR3[22] , \B_DOUT_TEMPR4[22] , \B_DOUT_TEMPR5[22] , 
        \B_DOUT_TEMPR6[22] , \B_DOUT_TEMPR7[22] , \B_DOUT_TEMPR8[22] , 
        \B_DOUT_TEMPR9[22] , \B_DOUT_TEMPR10[22] , 
        \B_DOUT_TEMPR11[22] , \B_DOUT_TEMPR12[22] , 
        \B_DOUT_TEMPR13[22] , \B_DOUT_TEMPR14[22] , 
        \B_DOUT_TEMPR15[22] , \B_DOUT_TEMPR16[22] , 
        \B_DOUT_TEMPR17[22] , \B_DOUT_TEMPR18[22] , 
        \B_DOUT_TEMPR19[22] , \B_DOUT_TEMPR20[22] , 
        \B_DOUT_TEMPR21[22] , \B_DOUT_TEMPR22[22] , 
        \B_DOUT_TEMPR23[22] , \B_DOUT_TEMPR24[22] , 
        \B_DOUT_TEMPR25[22] , \B_DOUT_TEMPR26[22] , 
        \B_DOUT_TEMPR27[22] , \B_DOUT_TEMPR28[22] , 
        \B_DOUT_TEMPR29[22] , \B_DOUT_TEMPR30[22] , 
        \B_DOUT_TEMPR31[22] , \B_DOUT_TEMPR32[22] , 
        \B_DOUT_TEMPR33[22] , \B_DOUT_TEMPR34[22] , 
        \B_DOUT_TEMPR35[22] , \B_DOUT_TEMPR36[22] , 
        \B_DOUT_TEMPR37[22] , \B_DOUT_TEMPR38[22] , 
        \B_DOUT_TEMPR39[22] , \B_DOUT_TEMPR40[22] , 
        \B_DOUT_TEMPR41[22] , \B_DOUT_TEMPR42[22] , 
        \B_DOUT_TEMPR43[22] , \B_DOUT_TEMPR44[22] , 
        \B_DOUT_TEMPR45[22] , \B_DOUT_TEMPR46[22] , 
        \B_DOUT_TEMPR47[22] , \B_DOUT_TEMPR48[22] , 
        \B_DOUT_TEMPR49[22] , \B_DOUT_TEMPR50[22] , 
        \B_DOUT_TEMPR51[22] , \B_DOUT_TEMPR52[22] , 
        \B_DOUT_TEMPR53[22] , \B_DOUT_TEMPR54[22] , 
        \B_DOUT_TEMPR55[22] , \B_DOUT_TEMPR56[22] , 
        \B_DOUT_TEMPR57[22] , \B_DOUT_TEMPR58[22] , 
        \B_DOUT_TEMPR59[22] , \B_DOUT_TEMPR60[22] , 
        \B_DOUT_TEMPR61[22] , \B_DOUT_TEMPR62[22] , 
        \B_DOUT_TEMPR63[22] , \B_DOUT_TEMPR64[22] , 
        \B_DOUT_TEMPR65[22] , \B_DOUT_TEMPR66[22] , 
        \B_DOUT_TEMPR67[22] , \B_DOUT_TEMPR68[22] , 
        \B_DOUT_TEMPR69[22] , \B_DOUT_TEMPR70[22] , 
        \B_DOUT_TEMPR71[22] , \B_DOUT_TEMPR72[22] , 
        \B_DOUT_TEMPR73[22] , \B_DOUT_TEMPR74[22] , 
        \B_DOUT_TEMPR75[22] , \B_DOUT_TEMPR76[22] , 
        \B_DOUT_TEMPR77[22] , \B_DOUT_TEMPR78[22] , 
        \B_DOUT_TEMPR79[22] , \B_DOUT_TEMPR80[22] , 
        \B_DOUT_TEMPR81[22] , \B_DOUT_TEMPR82[22] , 
        \B_DOUT_TEMPR83[22] , \B_DOUT_TEMPR84[22] , 
        \B_DOUT_TEMPR85[22] , \B_DOUT_TEMPR86[22] , 
        \B_DOUT_TEMPR87[22] , \B_DOUT_TEMPR88[22] , 
        \B_DOUT_TEMPR89[22] , \B_DOUT_TEMPR90[22] , 
        \B_DOUT_TEMPR91[22] , \B_DOUT_TEMPR92[22] , 
        \B_DOUT_TEMPR93[22] , \B_DOUT_TEMPR94[22] , 
        \B_DOUT_TEMPR95[22] , \B_DOUT_TEMPR96[22] , 
        \B_DOUT_TEMPR97[22] , \B_DOUT_TEMPR98[22] , 
        \B_DOUT_TEMPR99[22] , \B_DOUT_TEMPR100[22] , 
        \B_DOUT_TEMPR101[22] , \B_DOUT_TEMPR102[22] , 
        \B_DOUT_TEMPR103[22] , \B_DOUT_TEMPR104[22] , 
        \B_DOUT_TEMPR105[22] , \B_DOUT_TEMPR106[22] , 
        \B_DOUT_TEMPR107[22] , \B_DOUT_TEMPR108[22] , 
        \B_DOUT_TEMPR109[22] , \B_DOUT_TEMPR110[22] , 
        \B_DOUT_TEMPR111[22] , \B_DOUT_TEMPR112[22] , 
        \B_DOUT_TEMPR113[22] , \B_DOUT_TEMPR114[22] , 
        \B_DOUT_TEMPR115[22] , \B_DOUT_TEMPR116[22] , 
        \B_DOUT_TEMPR117[22] , \B_DOUT_TEMPR118[22] , 
        \B_DOUT_TEMPR0[23] , \B_DOUT_TEMPR1[23] , \B_DOUT_TEMPR2[23] , 
        \B_DOUT_TEMPR3[23] , \B_DOUT_TEMPR4[23] , \B_DOUT_TEMPR5[23] , 
        \B_DOUT_TEMPR6[23] , \B_DOUT_TEMPR7[23] , \B_DOUT_TEMPR8[23] , 
        \B_DOUT_TEMPR9[23] , \B_DOUT_TEMPR10[23] , 
        \B_DOUT_TEMPR11[23] , \B_DOUT_TEMPR12[23] , 
        \B_DOUT_TEMPR13[23] , \B_DOUT_TEMPR14[23] , 
        \B_DOUT_TEMPR15[23] , \B_DOUT_TEMPR16[23] , 
        \B_DOUT_TEMPR17[23] , \B_DOUT_TEMPR18[23] , 
        \B_DOUT_TEMPR19[23] , \B_DOUT_TEMPR20[23] , 
        \B_DOUT_TEMPR21[23] , \B_DOUT_TEMPR22[23] , 
        \B_DOUT_TEMPR23[23] , \B_DOUT_TEMPR24[23] , 
        \B_DOUT_TEMPR25[23] , \B_DOUT_TEMPR26[23] , 
        \B_DOUT_TEMPR27[23] , \B_DOUT_TEMPR28[23] , 
        \B_DOUT_TEMPR29[23] , \B_DOUT_TEMPR30[23] , 
        \B_DOUT_TEMPR31[23] , \B_DOUT_TEMPR32[23] , 
        \B_DOUT_TEMPR33[23] , \B_DOUT_TEMPR34[23] , 
        \B_DOUT_TEMPR35[23] , \B_DOUT_TEMPR36[23] , 
        \B_DOUT_TEMPR37[23] , \B_DOUT_TEMPR38[23] , 
        \B_DOUT_TEMPR39[23] , \B_DOUT_TEMPR40[23] , 
        \B_DOUT_TEMPR41[23] , \B_DOUT_TEMPR42[23] , 
        \B_DOUT_TEMPR43[23] , \B_DOUT_TEMPR44[23] , 
        \B_DOUT_TEMPR45[23] , \B_DOUT_TEMPR46[23] , 
        \B_DOUT_TEMPR47[23] , \B_DOUT_TEMPR48[23] , 
        \B_DOUT_TEMPR49[23] , \B_DOUT_TEMPR50[23] , 
        \B_DOUT_TEMPR51[23] , \B_DOUT_TEMPR52[23] , 
        \B_DOUT_TEMPR53[23] , \B_DOUT_TEMPR54[23] , 
        \B_DOUT_TEMPR55[23] , \B_DOUT_TEMPR56[23] , 
        \B_DOUT_TEMPR57[23] , \B_DOUT_TEMPR58[23] , 
        \B_DOUT_TEMPR59[23] , \B_DOUT_TEMPR60[23] , 
        \B_DOUT_TEMPR61[23] , \B_DOUT_TEMPR62[23] , 
        \B_DOUT_TEMPR63[23] , \B_DOUT_TEMPR64[23] , 
        \B_DOUT_TEMPR65[23] , \B_DOUT_TEMPR66[23] , 
        \B_DOUT_TEMPR67[23] , \B_DOUT_TEMPR68[23] , 
        \B_DOUT_TEMPR69[23] , \B_DOUT_TEMPR70[23] , 
        \B_DOUT_TEMPR71[23] , \B_DOUT_TEMPR72[23] , 
        \B_DOUT_TEMPR73[23] , \B_DOUT_TEMPR74[23] , 
        \B_DOUT_TEMPR75[23] , \B_DOUT_TEMPR76[23] , 
        \B_DOUT_TEMPR77[23] , \B_DOUT_TEMPR78[23] , 
        \B_DOUT_TEMPR79[23] , \B_DOUT_TEMPR80[23] , 
        \B_DOUT_TEMPR81[23] , \B_DOUT_TEMPR82[23] , 
        \B_DOUT_TEMPR83[23] , \B_DOUT_TEMPR84[23] , 
        \B_DOUT_TEMPR85[23] , \B_DOUT_TEMPR86[23] , 
        \B_DOUT_TEMPR87[23] , \B_DOUT_TEMPR88[23] , 
        \B_DOUT_TEMPR89[23] , \B_DOUT_TEMPR90[23] , 
        \B_DOUT_TEMPR91[23] , \B_DOUT_TEMPR92[23] , 
        \B_DOUT_TEMPR93[23] , \B_DOUT_TEMPR94[23] , 
        \B_DOUT_TEMPR95[23] , \B_DOUT_TEMPR96[23] , 
        \B_DOUT_TEMPR97[23] , \B_DOUT_TEMPR98[23] , 
        \B_DOUT_TEMPR99[23] , \B_DOUT_TEMPR100[23] , 
        \B_DOUT_TEMPR101[23] , \B_DOUT_TEMPR102[23] , 
        \B_DOUT_TEMPR103[23] , \B_DOUT_TEMPR104[23] , 
        \B_DOUT_TEMPR105[23] , \B_DOUT_TEMPR106[23] , 
        \B_DOUT_TEMPR107[23] , \B_DOUT_TEMPR108[23] , 
        \B_DOUT_TEMPR109[23] , \B_DOUT_TEMPR110[23] , 
        \B_DOUT_TEMPR111[23] , \B_DOUT_TEMPR112[23] , 
        \B_DOUT_TEMPR113[23] , \B_DOUT_TEMPR114[23] , 
        \B_DOUT_TEMPR115[23] , \B_DOUT_TEMPR116[23] , 
        \B_DOUT_TEMPR117[23] , \B_DOUT_TEMPR118[23] , 
        \B_DOUT_TEMPR0[24] , \B_DOUT_TEMPR1[24] , \B_DOUT_TEMPR2[24] , 
        \B_DOUT_TEMPR3[24] , \B_DOUT_TEMPR4[24] , \B_DOUT_TEMPR5[24] , 
        \B_DOUT_TEMPR6[24] , \B_DOUT_TEMPR7[24] , \B_DOUT_TEMPR8[24] , 
        \B_DOUT_TEMPR9[24] , \B_DOUT_TEMPR10[24] , 
        \B_DOUT_TEMPR11[24] , \B_DOUT_TEMPR12[24] , 
        \B_DOUT_TEMPR13[24] , \B_DOUT_TEMPR14[24] , 
        \B_DOUT_TEMPR15[24] , \B_DOUT_TEMPR16[24] , 
        \B_DOUT_TEMPR17[24] , \B_DOUT_TEMPR18[24] , 
        \B_DOUT_TEMPR19[24] , \B_DOUT_TEMPR20[24] , 
        \B_DOUT_TEMPR21[24] , \B_DOUT_TEMPR22[24] , 
        \B_DOUT_TEMPR23[24] , \B_DOUT_TEMPR24[24] , 
        \B_DOUT_TEMPR25[24] , \B_DOUT_TEMPR26[24] , 
        \B_DOUT_TEMPR27[24] , \B_DOUT_TEMPR28[24] , 
        \B_DOUT_TEMPR29[24] , \B_DOUT_TEMPR30[24] , 
        \B_DOUT_TEMPR31[24] , \B_DOUT_TEMPR32[24] , 
        \B_DOUT_TEMPR33[24] , \B_DOUT_TEMPR34[24] , 
        \B_DOUT_TEMPR35[24] , \B_DOUT_TEMPR36[24] , 
        \B_DOUT_TEMPR37[24] , \B_DOUT_TEMPR38[24] , 
        \B_DOUT_TEMPR39[24] , \B_DOUT_TEMPR40[24] , 
        \B_DOUT_TEMPR41[24] , \B_DOUT_TEMPR42[24] , 
        \B_DOUT_TEMPR43[24] , \B_DOUT_TEMPR44[24] , 
        \B_DOUT_TEMPR45[24] , \B_DOUT_TEMPR46[24] , 
        \B_DOUT_TEMPR47[24] , \B_DOUT_TEMPR48[24] , 
        \B_DOUT_TEMPR49[24] , \B_DOUT_TEMPR50[24] , 
        \B_DOUT_TEMPR51[24] , \B_DOUT_TEMPR52[24] , 
        \B_DOUT_TEMPR53[24] , \B_DOUT_TEMPR54[24] , 
        \B_DOUT_TEMPR55[24] , \B_DOUT_TEMPR56[24] , 
        \B_DOUT_TEMPR57[24] , \B_DOUT_TEMPR58[24] , 
        \B_DOUT_TEMPR59[24] , \B_DOUT_TEMPR60[24] , 
        \B_DOUT_TEMPR61[24] , \B_DOUT_TEMPR62[24] , 
        \B_DOUT_TEMPR63[24] , \B_DOUT_TEMPR64[24] , 
        \B_DOUT_TEMPR65[24] , \B_DOUT_TEMPR66[24] , 
        \B_DOUT_TEMPR67[24] , \B_DOUT_TEMPR68[24] , 
        \B_DOUT_TEMPR69[24] , \B_DOUT_TEMPR70[24] , 
        \B_DOUT_TEMPR71[24] , \B_DOUT_TEMPR72[24] , 
        \B_DOUT_TEMPR73[24] , \B_DOUT_TEMPR74[24] , 
        \B_DOUT_TEMPR75[24] , \B_DOUT_TEMPR76[24] , 
        \B_DOUT_TEMPR77[24] , \B_DOUT_TEMPR78[24] , 
        \B_DOUT_TEMPR79[24] , \B_DOUT_TEMPR80[24] , 
        \B_DOUT_TEMPR81[24] , \B_DOUT_TEMPR82[24] , 
        \B_DOUT_TEMPR83[24] , \B_DOUT_TEMPR84[24] , 
        \B_DOUT_TEMPR85[24] , \B_DOUT_TEMPR86[24] , 
        \B_DOUT_TEMPR87[24] , \B_DOUT_TEMPR88[24] , 
        \B_DOUT_TEMPR89[24] , \B_DOUT_TEMPR90[24] , 
        \B_DOUT_TEMPR91[24] , \B_DOUT_TEMPR92[24] , 
        \B_DOUT_TEMPR93[24] , \B_DOUT_TEMPR94[24] , 
        \B_DOUT_TEMPR95[24] , \B_DOUT_TEMPR96[24] , 
        \B_DOUT_TEMPR97[24] , \B_DOUT_TEMPR98[24] , 
        \B_DOUT_TEMPR99[24] , \B_DOUT_TEMPR100[24] , 
        \B_DOUT_TEMPR101[24] , \B_DOUT_TEMPR102[24] , 
        \B_DOUT_TEMPR103[24] , \B_DOUT_TEMPR104[24] , 
        \B_DOUT_TEMPR105[24] , \B_DOUT_TEMPR106[24] , 
        \B_DOUT_TEMPR107[24] , \B_DOUT_TEMPR108[24] , 
        \B_DOUT_TEMPR109[24] , \B_DOUT_TEMPR110[24] , 
        \B_DOUT_TEMPR111[24] , \B_DOUT_TEMPR112[24] , 
        \B_DOUT_TEMPR113[24] , \B_DOUT_TEMPR114[24] , 
        \B_DOUT_TEMPR115[24] , \B_DOUT_TEMPR116[24] , 
        \B_DOUT_TEMPR117[24] , \B_DOUT_TEMPR118[24] , 
        \B_DOUT_TEMPR0[25] , \B_DOUT_TEMPR1[25] , \B_DOUT_TEMPR2[25] , 
        \B_DOUT_TEMPR3[25] , \B_DOUT_TEMPR4[25] , \B_DOUT_TEMPR5[25] , 
        \B_DOUT_TEMPR6[25] , \B_DOUT_TEMPR7[25] , \B_DOUT_TEMPR8[25] , 
        \B_DOUT_TEMPR9[25] , \B_DOUT_TEMPR10[25] , 
        \B_DOUT_TEMPR11[25] , \B_DOUT_TEMPR12[25] , 
        \B_DOUT_TEMPR13[25] , \B_DOUT_TEMPR14[25] , 
        \B_DOUT_TEMPR15[25] , \B_DOUT_TEMPR16[25] , 
        \B_DOUT_TEMPR17[25] , \B_DOUT_TEMPR18[25] , 
        \B_DOUT_TEMPR19[25] , \B_DOUT_TEMPR20[25] , 
        \B_DOUT_TEMPR21[25] , \B_DOUT_TEMPR22[25] , 
        \B_DOUT_TEMPR23[25] , \B_DOUT_TEMPR24[25] , 
        \B_DOUT_TEMPR25[25] , \B_DOUT_TEMPR26[25] , 
        \B_DOUT_TEMPR27[25] , \B_DOUT_TEMPR28[25] , 
        \B_DOUT_TEMPR29[25] , \B_DOUT_TEMPR30[25] , 
        \B_DOUT_TEMPR31[25] , \B_DOUT_TEMPR32[25] , 
        \B_DOUT_TEMPR33[25] , \B_DOUT_TEMPR34[25] , 
        \B_DOUT_TEMPR35[25] , \B_DOUT_TEMPR36[25] , 
        \B_DOUT_TEMPR37[25] , \B_DOUT_TEMPR38[25] , 
        \B_DOUT_TEMPR39[25] , \B_DOUT_TEMPR40[25] , 
        \B_DOUT_TEMPR41[25] , \B_DOUT_TEMPR42[25] , 
        \B_DOUT_TEMPR43[25] , \B_DOUT_TEMPR44[25] , 
        \B_DOUT_TEMPR45[25] , \B_DOUT_TEMPR46[25] , 
        \B_DOUT_TEMPR47[25] , \B_DOUT_TEMPR48[25] , 
        \B_DOUT_TEMPR49[25] , \B_DOUT_TEMPR50[25] , 
        \B_DOUT_TEMPR51[25] , \B_DOUT_TEMPR52[25] , 
        \B_DOUT_TEMPR53[25] , \B_DOUT_TEMPR54[25] , 
        \B_DOUT_TEMPR55[25] , \B_DOUT_TEMPR56[25] , 
        \B_DOUT_TEMPR57[25] , \B_DOUT_TEMPR58[25] , 
        \B_DOUT_TEMPR59[25] , \B_DOUT_TEMPR60[25] , 
        \B_DOUT_TEMPR61[25] , \B_DOUT_TEMPR62[25] , 
        \B_DOUT_TEMPR63[25] , \B_DOUT_TEMPR64[25] , 
        \B_DOUT_TEMPR65[25] , \B_DOUT_TEMPR66[25] , 
        \B_DOUT_TEMPR67[25] , \B_DOUT_TEMPR68[25] , 
        \B_DOUT_TEMPR69[25] , \B_DOUT_TEMPR70[25] , 
        \B_DOUT_TEMPR71[25] , \B_DOUT_TEMPR72[25] , 
        \B_DOUT_TEMPR73[25] , \B_DOUT_TEMPR74[25] , 
        \B_DOUT_TEMPR75[25] , \B_DOUT_TEMPR76[25] , 
        \B_DOUT_TEMPR77[25] , \B_DOUT_TEMPR78[25] , 
        \B_DOUT_TEMPR79[25] , \B_DOUT_TEMPR80[25] , 
        \B_DOUT_TEMPR81[25] , \B_DOUT_TEMPR82[25] , 
        \B_DOUT_TEMPR83[25] , \B_DOUT_TEMPR84[25] , 
        \B_DOUT_TEMPR85[25] , \B_DOUT_TEMPR86[25] , 
        \B_DOUT_TEMPR87[25] , \B_DOUT_TEMPR88[25] , 
        \B_DOUT_TEMPR89[25] , \B_DOUT_TEMPR90[25] , 
        \B_DOUT_TEMPR91[25] , \B_DOUT_TEMPR92[25] , 
        \B_DOUT_TEMPR93[25] , \B_DOUT_TEMPR94[25] , 
        \B_DOUT_TEMPR95[25] , \B_DOUT_TEMPR96[25] , 
        \B_DOUT_TEMPR97[25] , \B_DOUT_TEMPR98[25] , 
        \B_DOUT_TEMPR99[25] , \B_DOUT_TEMPR100[25] , 
        \B_DOUT_TEMPR101[25] , \B_DOUT_TEMPR102[25] , 
        \B_DOUT_TEMPR103[25] , \B_DOUT_TEMPR104[25] , 
        \B_DOUT_TEMPR105[25] , \B_DOUT_TEMPR106[25] , 
        \B_DOUT_TEMPR107[25] , \B_DOUT_TEMPR108[25] , 
        \B_DOUT_TEMPR109[25] , \B_DOUT_TEMPR110[25] , 
        \B_DOUT_TEMPR111[25] , \B_DOUT_TEMPR112[25] , 
        \B_DOUT_TEMPR113[25] , \B_DOUT_TEMPR114[25] , 
        \B_DOUT_TEMPR115[25] , \B_DOUT_TEMPR116[25] , 
        \B_DOUT_TEMPR117[25] , \B_DOUT_TEMPR118[25] , 
        \B_DOUT_TEMPR0[26] , \B_DOUT_TEMPR1[26] , \B_DOUT_TEMPR2[26] , 
        \B_DOUT_TEMPR3[26] , \B_DOUT_TEMPR4[26] , \B_DOUT_TEMPR5[26] , 
        \B_DOUT_TEMPR6[26] , \B_DOUT_TEMPR7[26] , \B_DOUT_TEMPR8[26] , 
        \B_DOUT_TEMPR9[26] , \B_DOUT_TEMPR10[26] , 
        \B_DOUT_TEMPR11[26] , \B_DOUT_TEMPR12[26] , 
        \B_DOUT_TEMPR13[26] , \B_DOUT_TEMPR14[26] , 
        \B_DOUT_TEMPR15[26] , \B_DOUT_TEMPR16[26] , 
        \B_DOUT_TEMPR17[26] , \B_DOUT_TEMPR18[26] , 
        \B_DOUT_TEMPR19[26] , \B_DOUT_TEMPR20[26] , 
        \B_DOUT_TEMPR21[26] , \B_DOUT_TEMPR22[26] , 
        \B_DOUT_TEMPR23[26] , \B_DOUT_TEMPR24[26] , 
        \B_DOUT_TEMPR25[26] , \B_DOUT_TEMPR26[26] , 
        \B_DOUT_TEMPR27[26] , \B_DOUT_TEMPR28[26] , 
        \B_DOUT_TEMPR29[26] , \B_DOUT_TEMPR30[26] , 
        \B_DOUT_TEMPR31[26] , \B_DOUT_TEMPR32[26] , 
        \B_DOUT_TEMPR33[26] , \B_DOUT_TEMPR34[26] , 
        \B_DOUT_TEMPR35[26] , \B_DOUT_TEMPR36[26] , 
        \B_DOUT_TEMPR37[26] , \B_DOUT_TEMPR38[26] , 
        \B_DOUT_TEMPR39[26] , \B_DOUT_TEMPR40[26] , 
        \B_DOUT_TEMPR41[26] , \B_DOUT_TEMPR42[26] , 
        \B_DOUT_TEMPR43[26] , \B_DOUT_TEMPR44[26] , 
        \B_DOUT_TEMPR45[26] , \B_DOUT_TEMPR46[26] , 
        \B_DOUT_TEMPR47[26] , \B_DOUT_TEMPR48[26] , 
        \B_DOUT_TEMPR49[26] , \B_DOUT_TEMPR50[26] , 
        \B_DOUT_TEMPR51[26] , \B_DOUT_TEMPR52[26] , 
        \B_DOUT_TEMPR53[26] , \B_DOUT_TEMPR54[26] , 
        \B_DOUT_TEMPR55[26] , \B_DOUT_TEMPR56[26] , 
        \B_DOUT_TEMPR57[26] , \B_DOUT_TEMPR58[26] , 
        \B_DOUT_TEMPR59[26] , \B_DOUT_TEMPR60[26] , 
        \B_DOUT_TEMPR61[26] , \B_DOUT_TEMPR62[26] , 
        \B_DOUT_TEMPR63[26] , \B_DOUT_TEMPR64[26] , 
        \B_DOUT_TEMPR65[26] , \B_DOUT_TEMPR66[26] , 
        \B_DOUT_TEMPR67[26] , \B_DOUT_TEMPR68[26] , 
        \B_DOUT_TEMPR69[26] , \B_DOUT_TEMPR70[26] , 
        \B_DOUT_TEMPR71[26] , \B_DOUT_TEMPR72[26] , 
        \B_DOUT_TEMPR73[26] , \B_DOUT_TEMPR74[26] , 
        \B_DOUT_TEMPR75[26] , \B_DOUT_TEMPR76[26] , 
        \B_DOUT_TEMPR77[26] , \B_DOUT_TEMPR78[26] , 
        \B_DOUT_TEMPR79[26] , \B_DOUT_TEMPR80[26] , 
        \B_DOUT_TEMPR81[26] , \B_DOUT_TEMPR82[26] , 
        \B_DOUT_TEMPR83[26] , \B_DOUT_TEMPR84[26] , 
        \B_DOUT_TEMPR85[26] , \B_DOUT_TEMPR86[26] , 
        \B_DOUT_TEMPR87[26] , \B_DOUT_TEMPR88[26] , 
        \B_DOUT_TEMPR89[26] , \B_DOUT_TEMPR90[26] , 
        \B_DOUT_TEMPR91[26] , \B_DOUT_TEMPR92[26] , 
        \B_DOUT_TEMPR93[26] , \B_DOUT_TEMPR94[26] , 
        \B_DOUT_TEMPR95[26] , \B_DOUT_TEMPR96[26] , 
        \B_DOUT_TEMPR97[26] , \B_DOUT_TEMPR98[26] , 
        \B_DOUT_TEMPR99[26] , \B_DOUT_TEMPR100[26] , 
        \B_DOUT_TEMPR101[26] , \B_DOUT_TEMPR102[26] , 
        \B_DOUT_TEMPR103[26] , \B_DOUT_TEMPR104[26] , 
        \B_DOUT_TEMPR105[26] , \B_DOUT_TEMPR106[26] , 
        \B_DOUT_TEMPR107[26] , \B_DOUT_TEMPR108[26] , 
        \B_DOUT_TEMPR109[26] , \B_DOUT_TEMPR110[26] , 
        \B_DOUT_TEMPR111[26] , \B_DOUT_TEMPR112[26] , 
        \B_DOUT_TEMPR113[26] , \B_DOUT_TEMPR114[26] , 
        \B_DOUT_TEMPR115[26] , \B_DOUT_TEMPR116[26] , 
        \B_DOUT_TEMPR117[26] , \B_DOUT_TEMPR118[26] , 
        \B_DOUT_TEMPR0[27] , \B_DOUT_TEMPR1[27] , \B_DOUT_TEMPR2[27] , 
        \B_DOUT_TEMPR3[27] , \B_DOUT_TEMPR4[27] , \B_DOUT_TEMPR5[27] , 
        \B_DOUT_TEMPR6[27] , \B_DOUT_TEMPR7[27] , \B_DOUT_TEMPR8[27] , 
        \B_DOUT_TEMPR9[27] , \B_DOUT_TEMPR10[27] , 
        \B_DOUT_TEMPR11[27] , \B_DOUT_TEMPR12[27] , 
        \B_DOUT_TEMPR13[27] , \B_DOUT_TEMPR14[27] , 
        \B_DOUT_TEMPR15[27] , \B_DOUT_TEMPR16[27] , 
        \B_DOUT_TEMPR17[27] , \B_DOUT_TEMPR18[27] , 
        \B_DOUT_TEMPR19[27] , \B_DOUT_TEMPR20[27] , 
        \B_DOUT_TEMPR21[27] , \B_DOUT_TEMPR22[27] , 
        \B_DOUT_TEMPR23[27] , \B_DOUT_TEMPR24[27] , 
        \B_DOUT_TEMPR25[27] , \B_DOUT_TEMPR26[27] , 
        \B_DOUT_TEMPR27[27] , \B_DOUT_TEMPR28[27] , 
        \B_DOUT_TEMPR29[27] , \B_DOUT_TEMPR30[27] , 
        \B_DOUT_TEMPR31[27] , \B_DOUT_TEMPR32[27] , 
        \B_DOUT_TEMPR33[27] , \B_DOUT_TEMPR34[27] , 
        \B_DOUT_TEMPR35[27] , \B_DOUT_TEMPR36[27] , 
        \B_DOUT_TEMPR37[27] , \B_DOUT_TEMPR38[27] , 
        \B_DOUT_TEMPR39[27] , \B_DOUT_TEMPR40[27] , 
        \B_DOUT_TEMPR41[27] , \B_DOUT_TEMPR42[27] , 
        \B_DOUT_TEMPR43[27] , \B_DOUT_TEMPR44[27] , 
        \B_DOUT_TEMPR45[27] , \B_DOUT_TEMPR46[27] , 
        \B_DOUT_TEMPR47[27] , \B_DOUT_TEMPR48[27] , 
        \B_DOUT_TEMPR49[27] , \B_DOUT_TEMPR50[27] , 
        \B_DOUT_TEMPR51[27] , \B_DOUT_TEMPR52[27] , 
        \B_DOUT_TEMPR53[27] , \B_DOUT_TEMPR54[27] , 
        \B_DOUT_TEMPR55[27] , \B_DOUT_TEMPR56[27] , 
        \B_DOUT_TEMPR57[27] , \B_DOUT_TEMPR58[27] , 
        \B_DOUT_TEMPR59[27] , \B_DOUT_TEMPR60[27] , 
        \B_DOUT_TEMPR61[27] , \B_DOUT_TEMPR62[27] , 
        \B_DOUT_TEMPR63[27] , \B_DOUT_TEMPR64[27] , 
        \B_DOUT_TEMPR65[27] , \B_DOUT_TEMPR66[27] , 
        \B_DOUT_TEMPR67[27] , \B_DOUT_TEMPR68[27] , 
        \B_DOUT_TEMPR69[27] , \B_DOUT_TEMPR70[27] , 
        \B_DOUT_TEMPR71[27] , \B_DOUT_TEMPR72[27] , 
        \B_DOUT_TEMPR73[27] , \B_DOUT_TEMPR74[27] , 
        \B_DOUT_TEMPR75[27] , \B_DOUT_TEMPR76[27] , 
        \B_DOUT_TEMPR77[27] , \B_DOUT_TEMPR78[27] , 
        \B_DOUT_TEMPR79[27] , \B_DOUT_TEMPR80[27] , 
        \B_DOUT_TEMPR81[27] , \B_DOUT_TEMPR82[27] , 
        \B_DOUT_TEMPR83[27] , \B_DOUT_TEMPR84[27] , 
        \B_DOUT_TEMPR85[27] , \B_DOUT_TEMPR86[27] , 
        \B_DOUT_TEMPR87[27] , \B_DOUT_TEMPR88[27] , 
        \B_DOUT_TEMPR89[27] , \B_DOUT_TEMPR90[27] , 
        \B_DOUT_TEMPR91[27] , \B_DOUT_TEMPR92[27] , 
        \B_DOUT_TEMPR93[27] , \B_DOUT_TEMPR94[27] , 
        \B_DOUT_TEMPR95[27] , \B_DOUT_TEMPR96[27] , 
        \B_DOUT_TEMPR97[27] , \B_DOUT_TEMPR98[27] , 
        \B_DOUT_TEMPR99[27] , \B_DOUT_TEMPR100[27] , 
        \B_DOUT_TEMPR101[27] , \B_DOUT_TEMPR102[27] , 
        \B_DOUT_TEMPR103[27] , \B_DOUT_TEMPR104[27] , 
        \B_DOUT_TEMPR105[27] , \B_DOUT_TEMPR106[27] , 
        \B_DOUT_TEMPR107[27] , \B_DOUT_TEMPR108[27] , 
        \B_DOUT_TEMPR109[27] , \B_DOUT_TEMPR110[27] , 
        \B_DOUT_TEMPR111[27] , \B_DOUT_TEMPR112[27] , 
        \B_DOUT_TEMPR113[27] , \B_DOUT_TEMPR114[27] , 
        \B_DOUT_TEMPR115[27] , \B_DOUT_TEMPR116[27] , 
        \B_DOUT_TEMPR117[27] , \B_DOUT_TEMPR118[27] , 
        \B_DOUT_TEMPR0[28] , \B_DOUT_TEMPR1[28] , \B_DOUT_TEMPR2[28] , 
        \B_DOUT_TEMPR3[28] , \B_DOUT_TEMPR4[28] , \B_DOUT_TEMPR5[28] , 
        \B_DOUT_TEMPR6[28] , \B_DOUT_TEMPR7[28] , \B_DOUT_TEMPR8[28] , 
        \B_DOUT_TEMPR9[28] , \B_DOUT_TEMPR10[28] , 
        \B_DOUT_TEMPR11[28] , \B_DOUT_TEMPR12[28] , 
        \B_DOUT_TEMPR13[28] , \B_DOUT_TEMPR14[28] , 
        \B_DOUT_TEMPR15[28] , \B_DOUT_TEMPR16[28] , 
        \B_DOUT_TEMPR17[28] , \B_DOUT_TEMPR18[28] , 
        \B_DOUT_TEMPR19[28] , \B_DOUT_TEMPR20[28] , 
        \B_DOUT_TEMPR21[28] , \B_DOUT_TEMPR22[28] , 
        \B_DOUT_TEMPR23[28] , \B_DOUT_TEMPR24[28] , 
        \B_DOUT_TEMPR25[28] , \B_DOUT_TEMPR26[28] , 
        \B_DOUT_TEMPR27[28] , \B_DOUT_TEMPR28[28] , 
        \B_DOUT_TEMPR29[28] , \B_DOUT_TEMPR30[28] , 
        \B_DOUT_TEMPR31[28] , \B_DOUT_TEMPR32[28] , 
        \B_DOUT_TEMPR33[28] , \B_DOUT_TEMPR34[28] , 
        \B_DOUT_TEMPR35[28] , \B_DOUT_TEMPR36[28] , 
        \B_DOUT_TEMPR37[28] , \B_DOUT_TEMPR38[28] , 
        \B_DOUT_TEMPR39[28] , \B_DOUT_TEMPR40[28] , 
        \B_DOUT_TEMPR41[28] , \B_DOUT_TEMPR42[28] , 
        \B_DOUT_TEMPR43[28] , \B_DOUT_TEMPR44[28] , 
        \B_DOUT_TEMPR45[28] , \B_DOUT_TEMPR46[28] , 
        \B_DOUT_TEMPR47[28] , \B_DOUT_TEMPR48[28] , 
        \B_DOUT_TEMPR49[28] , \B_DOUT_TEMPR50[28] , 
        \B_DOUT_TEMPR51[28] , \B_DOUT_TEMPR52[28] , 
        \B_DOUT_TEMPR53[28] , \B_DOUT_TEMPR54[28] , 
        \B_DOUT_TEMPR55[28] , \B_DOUT_TEMPR56[28] , 
        \B_DOUT_TEMPR57[28] , \B_DOUT_TEMPR58[28] , 
        \B_DOUT_TEMPR59[28] , \B_DOUT_TEMPR60[28] , 
        \B_DOUT_TEMPR61[28] , \B_DOUT_TEMPR62[28] , 
        \B_DOUT_TEMPR63[28] , \B_DOUT_TEMPR64[28] , 
        \B_DOUT_TEMPR65[28] , \B_DOUT_TEMPR66[28] , 
        \B_DOUT_TEMPR67[28] , \B_DOUT_TEMPR68[28] , 
        \B_DOUT_TEMPR69[28] , \B_DOUT_TEMPR70[28] , 
        \B_DOUT_TEMPR71[28] , \B_DOUT_TEMPR72[28] , 
        \B_DOUT_TEMPR73[28] , \B_DOUT_TEMPR74[28] , 
        \B_DOUT_TEMPR75[28] , \B_DOUT_TEMPR76[28] , 
        \B_DOUT_TEMPR77[28] , \B_DOUT_TEMPR78[28] , 
        \B_DOUT_TEMPR79[28] , \B_DOUT_TEMPR80[28] , 
        \B_DOUT_TEMPR81[28] , \B_DOUT_TEMPR82[28] , 
        \B_DOUT_TEMPR83[28] , \B_DOUT_TEMPR84[28] , 
        \B_DOUT_TEMPR85[28] , \B_DOUT_TEMPR86[28] , 
        \B_DOUT_TEMPR87[28] , \B_DOUT_TEMPR88[28] , 
        \B_DOUT_TEMPR89[28] , \B_DOUT_TEMPR90[28] , 
        \B_DOUT_TEMPR91[28] , \B_DOUT_TEMPR92[28] , 
        \B_DOUT_TEMPR93[28] , \B_DOUT_TEMPR94[28] , 
        \B_DOUT_TEMPR95[28] , \B_DOUT_TEMPR96[28] , 
        \B_DOUT_TEMPR97[28] , \B_DOUT_TEMPR98[28] , 
        \B_DOUT_TEMPR99[28] , \B_DOUT_TEMPR100[28] , 
        \B_DOUT_TEMPR101[28] , \B_DOUT_TEMPR102[28] , 
        \B_DOUT_TEMPR103[28] , \B_DOUT_TEMPR104[28] , 
        \B_DOUT_TEMPR105[28] , \B_DOUT_TEMPR106[28] , 
        \B_DOUT_TEMPR107[28] , \B_DOUT_TEMPR108[28] , 
        \B_DOUT_TEMPR109[28] , \B_DOUT_TEMPR110[28] , 
        \B_DOUT_TEMPR111[28] , \B_DOUT_TEMPR112[28] , 
        \B_DOUT_TEMPR113[28] , \B_DOUT_TEMPR114[28] , 
        \B_DOUT_TEMPR115[28] , \B_DOUT_TEMPR116[28] , 
        \B_DOUT_TEMPR117[28] , \B_DOUT_TEMPR118[28] , 
        \B_DOUT_TEMPR0[29] , \B_DOUT_TEMPR1[29] , \B_DOUT_TEMPR2[29] , 
        \B_DOUT_TEMPR3[29] , \B_DOUT_TEMPR4[29] , \B_DOUT_TEMPR5[29] , 
        \B_DOUT_TEMPR6[29] , \B_DOUT_TEMPR7[29] , \B_DOUT_TEMPR8[29] , 
        \B_DOUT_TEMPR9[29] , \B_DOUT_TEMPR10[29] , 
        \B_DOUT_TEMPR11[29] , \B_DOUT_TEMPR12[29] , 
        \B_DOUT_TEMPR13[29] , \B_DOUT_TEMPR14[29] , 
        \B_DOUT_TEMPR15[29] , \B_DOUT_TEMPR16[29] , 
        \B_DOUT_TEMPR17[29] , \B_DOUT_TEMPR18[29] , 
        \B_DOUT_TEMPR19[29] , \B_DOUT_TEMPR20[29] , 
        \B_DOUT_TEMPR21[29] , \B_DOUT_TEMPR22[29] , 
        \B_DOUT_TEMPR23[29] , \B_DOUT_TEMPR24[29] , 
        \B_DOUT_TEMPR25[29] , \B_DOUT_TEMPR26[29] , 
        \B_DOUT_TEMPR27[29] , \B_DOUT_TEMPR28[29] , 
        \B_DOUT_TEMPR29[29] , \B_DOUT_TEMPR30[29] , 
        \B_DOUT_TEMPR31[29] , \B_DOUT_TEMPR32[29] , 
        \B_DOUT_TEMPR33[29] , \B_DOUT_TEMPR34[29] , 
        \B_DOUT_TEMPR35[29] , \B_DOUT_TEMPR36[29] , 
        \B_DOUT_TEMPR37[29] , \B_DOUT_TEMPR38[29] , 
        \B_DOUT_TEMPR39[29] , \B_DOUT_TEMPR40[29] , 
        \B_DOUT_TEMPR41[29] , \B_DOUT_TEMPR42[29] , 
        \B_DOUT_TEMPR43[29] , \B_DOUT_TEMPR44[29] , 
        \B_DOUT_TEMPR45[29] , \B_DOUT_TEMPR46[29] , 
        \B_DOUT_TEMPR47[29] , \B_DOUT_TEMPR48[29] , 
        \B_DOUT_TEMPR49[29] , \B_DOUT_TEMPR50[29] , 
        \B_DOUT_TEMPR51[29] , \B_DOUT_TEMPR52[29] , 
        \B_DOUT_TEMPR53[29] , \B_DOUT_TEMPR54[29] , 
        \B_DOUT_TEMPR55[29] , \B_DOUT_TEMPR56[29] , 
        \B_DOUT_TEMPR57[29] , \B_DOUT_TEMPR58[29] , 
        \B_DOUT_TEMPR59[29] , \B_DOUT_TEMPR60[29] , 
        \B_DOUT_TEMPR61[29] , \B_DOUT_TEMPR62[29] , 
        \B_DOUT_TEMPR63[29] , \B_DOUT_TEMPR64[29] , 
        \B_DOUT_TEMPR65[29] , \B_DOUT_TEMPR66[29] , 
        \B_DOUT_TEMPR67[29] , \B_DOUT_TEMPR68[29] , 
        \B_DOUT_TEMPR69[29] , \B_DOUT_TEMPR70[29] , 
        \B_DOUT_TEMPR71[29] , \B_DOUT_TEMPR72[29] , 
        \B_DOUT_TEMPR73[29] , \B_DOUT_TEMPR74[29] , 
        \B_DOUT_TEMPR75[29] , \B_DOUT_TEMPR76[29] , 
        \B_DOUT_TEMPR77[29] , \B_DOUT_TEMPR78[29] , 
        \B_DOUT_TEMPR79[29] , \B_DOUT_TEMPR80[29] , 
        \B_DOUT_TEMPR81[29] , \B_DOUT_TEMPR82[29] , 
        \B_DOUT_TEMPR83[29] , \B_DOUT_TEMPR84[29] , 
        \B_DOUT_TEMPR85[29] , \B_DOUT_TEMPR86[29] , 
        \B_DOUT_TEMPR87[29] , \B_DOUT_TEMPR88[29] , 
        \B_DOUT_TEMPR89[29] , \B_DOUT_TEMPR90[29] , 
        \B_DOUT_TEMPR91[29] , \B_DOUT_TEMPR92[29] , 
        \B_DOUT_TEMPR93[29] , \B_DOUT_TEMPR94[29] , 
        \B_DOUT_TEMPR95[29] , \B_DOUT_TEMPR96[29] , 
        \B_DOUT_TEMPR97[29] , \B_DOUT_TEMPR98[29] , 
        \B_DOUT_TEMPR99[29] , \B_DOUT_TEMPR100[29] , 
        \B_DOUT_TEMPR101[29] , \B_DOUT_TEMPR102[29] , 
        \B_DOUT_TEMPR103[29] , \B_DOUT_TEMPR104[29] , 
        \B_DOUT_TEMPR105[29] , \B_DOUT_TEMPR106[29] , 
        \B_DOUT_TEMPR107[29] , \B_DOUT_TEMPR108[29] , 
        \B_DOUT_TEMPR109[29] , \B_DOUT_TEMPR110[29] , 
        \B_DOUT_TEMPR111[29] , \B_DOUT_TEMPR112[29] , 
        \B_DOUT_TEMPR113[29] , \B_DOUT_TEMPR114[29] , 
        \B_DOUT_TEMPR115[29] , \B_DOUT_TEMPR116[29] , 
        \B_DOUT_TEMPR117[29] , \B_DOUT_TEMPR118[29] , 
        \B_DOUT_TEMPR0[30] , \B_DOUT_TEMPR1[30] , \B_DOUT_TEMPR2[30] , 
        \B_DOUT_TEMPR3[30] , \B_DOUT_TEMPR4[30] , \B_DOUT_TEMPR5[30] , 
        \B_DOUT_TEMPR6[30] , \B_DOUT_TEMPR7[30] , \B_DOUT_TEMPR8[30] , 
        \B_DOUT_TEMPR9[30] , \B_DOUT_TEMPR10[30] , 
        \B_DOUT_TEMPR11[30] , \B_DOUT_TEMPR12[30] , 
        \B_DOUT_TEMPR13[30] , \B_DOUT_TEMPR14[30] , 
        \B_DOUT_TEMPR15[30] , \B_DOUT_TEMPR16[30] , 
        \B_DOUT_TEMPR17[30] , \B_DOUT_TEMPR18[30] , 
        \B_DOUT_TEMPR19[30] , \B_DOUT_TEMPR20[30] , 
        \B_DOUT_TEMPR21[30] , \B_DOUT_TEMPR22[30] , 
        \B_DOUT_TEMPR23[30] , \B_DOUT_TEMPR24[30] , 
        \B_DOUT_TEMPR25[30] , \B_DOUT_TEMPR26[30] , 
        \B_DOUT_TEMPR27[30] , \B_DOUT_TEMPR28[30] , 
        \B_DOUT_TEMPR29[30] , \B_DOUT_TEMPR30[30] , 
        \B_DOUT_TEMPR31[30] , \B_DOUT_TEMPR32[30] , 
        \B_DOUT_TEMPR33[30] , \B_DOUT_TEMPR34[30] , 
        \B_DOUT_TEMPR35[30] , \B_DOUT_TEMPR36[30] , 
        \B_DOUT_TEMPR37[30] , \B_DOUT_TEMPR38[30] , 
        \B_DOUT_TEMPR39[30] , \B_DOUT_TEMPR40[30] , 
        \B_DOUT_TEMPR41[30] , \B_DOUT_TEMPR42[30] , 
        \B_DOUT_TEMPR43[30] , \B_DOUT_TEMPR44[30] , 
        \B_DOUT_TEMPR45[30] , \B_DOUT_TEMPR46[30] , 
        \B_DOUT_TEMPR47[30] , \B_DOUT_TEMPR48[30] , 
        \B_DOUT_TEMPR49[30] , \B_DOUT_TEMPR50[30] , 
        \B_DOUT_TEMPR51[30] , \B_DOUT_TEMPR52[30] , 
        \B_DOUT_TEMPR53[30] , \B_DOUT_TEMPR54[30] , 
        \B_DOUT_TEMPR55[30] , \B_DOUT_TEMPR56[30] , 
        \B_DOUT_TEMPR57[30] , \B_DOUT_TEMPR58[30] , 
        \B_DOUT_TEMPR59[30] , \B_DOUT_TEMPR60[30] , 
        \B_DOUT_TEMPR61[30] , \B_DOUT_TEMPR62[30] , 
        \B_DOUT_TEMPR63[30] , \B_DOUT_TEMPR64[30] , 
        \B_DOUT_TEMPR65[30] , \B_DOUT_TEMPR66[30] , 
        \B_DOUT_TEMPR67[30] , \B_DOUT_TEMPR68[30] , 
        \B_DOUT_TEMPR69[30] , \B_DOUT_TEMPR70[30] , 
        \B_DOUT_TEMPR71[30] , \B_DOUT_TEMPR72[30] , 
        \B_DOUT_TEMPR73[30] , \B_DOUT_TEMPR74[30] , 
        \B_DOUT_TEMPR75[30] , \B_DOUT_TEMPR76[30] , 
        \B_DOUT_TEMPR77[30] , \B_DOUT_TEMPR78[30] , 
        \B_DOUT_TEMPR79[30] , \B_DOUT_TEMPR80[30] , 
        \B_DOUT_TEMPR81[30] , \B_DOUT_TEMPR82[30] , 
        \B_DOUT_TEMPR83[30] , \B_DOUT_TEMPR84[30] , 
        \B_DOUT_TEMPR85[30] , \B_DOUT_TEMPR86[30] , 
        \B_DOUT_TEMPR87[30] , \B_DOUT_TEMPR88[30] , 
        \B_DOUT_TEMPR89[30] , \B_DOUT_TEMPR90[30] , 
        \B_DOUT_TEMPR91[30] , \B_DOUT_TEMPR92[30] , 
        \B_DOUT_TEMPR93[30] , \B_DOUT_TEMPR94[30] , 
        \B_DOUT_TEMPR95[30] , \B_DOUT_TEMPR96[30] , 
        \B_DOUT_TEMPR97[30] , \B_DOUT_TEMPR98[30] , 
        \B_DOUT_TEMPR99[30] , \B_DOUT_TEMPR100[30] , 
        \B_DOUT_TEMPR101[30] , \B_DOUT_TEMPR102[30] , 
        \B_DOUT_TEMPR103[30] , \B_DOUT_TEMPR104[30] , 
        \B_DOUT_TEMPR105[30] , \B_DOUT_TEMPR106[30] , 
        \B_DOUT_TEMPR107[30] , \B_DOUT_TEMPR108[30] , 
        \B_DOUT_TEMPR109[30] , \B_DOUT_TEMPR110[30] , 
        \B_DOUT_TEMPR111[30] , \B_DOUT_TEMPR112[30] , 
        \B_DOUT_TEMPR113[30] , \B_DOUT_TEMPR114[30] , 
        \B_DOUT_TEMPR115[30] , \B_DOUT_TEMPR116[30] , 
        \B_DOUT_TEMPR117[30] , \B_DOUT_TEMPR118[30] , 
        \B_DOUT_TEMPR0[31] , \B_DOUT_TEMPR1[31] , \B_DOUT_TEMPR2[31] , 
        \B_DOUT_TEMPR3[31] , \B_DOUT_TEMPR4[31] , \B_DOUT_TEMPR5[31] , 
        \B_DOUT_TEMPR6[31] , \B_DOUT_TEMPR7[31] , \B_DOUT_TEMPR8[31] , 
        \B_DOUT_TEMPR9[31] , \B_DOUT_TEMPR10[31] , 
        \B_DOUT_TEMPR11[31] , \B_DOUT_TEMPR12[31] , 
        \B_DOUT_TEMPR13[31] , \B_DOUT_TEMPR14[31] , 
        \B_DOUT_TEMPR15[31] , \B_DOUT_TEMPR16[31] , 
        \B_DOUT_TEMPR17[31] , \B_DOUT_TEMPR18[31] , 
        \B_DOUT_TEMPR19[31] , \B_DOUT_TEMPR20[31] , 
        \B_DOUT_TEMPR21[31] , \B_DOUT_TEMPR22[31] , 
        \B_DOUT_TEMPR23[31] , \B_DOUT_TEMPR24[31] , 
        \B_DOUT_TEMPR25[31] , \B_DOUT_TEMPR26[31] , 
        \B_DOUT_TEMPR27[31] , \B_DOUT_TEMPR28[31] , 
        \B_DOUT_TEMPR29[31] , \B_DOUT_TEMPR30[31] , 
        \B_DOUT_TEMPR31[31] , \B_DOUT_TEMPR32[31] , 
        \B_DOUT_TEMPR33[31] , \B_DOUT_TEMPR34[31] , 
        \B_DOUT_TEMPR35[31] , \B_DOUT_TEMPR36[31] , 
        \B_DOUT_TEMPR37[31] , \B_DOUT_TEMPR38[31] , 
        \B_DOUT_TEMPR39[31] , \B_DOUT_TEMPR40[31] , 
        \B_DOUT_TEMPR41[31] , \B_DOUT_TEMPR42[31] , 
        \B_DOUT_TEMPR43[31] , \B_DOUT_TEMPR44[31] , 
        \B_DOUT_TEMPR45[31] , \B_DOUT_TEMPR46[31] , 
        \B_DOUT_TEMPR47[31] , \B_DOUT_TEMPR48[31] , 
        \B_DOUT_TEMPR49[31] , \B_DOUT_TEMPR50[31] , 
        \B_DOUT_TEMPR51[31] , \B_DOUT_TEMPR52[31] , 
        \B_DOUT_TEMPR53[31] , \B_DOUT_TEMPR54[31] , 
        \B_DOUT_TEMPR55[31] , \B_DOUT_TEMPR56[31] , 
        \B_DOUT_TEMPR57[31] , \B_DOUT_TEMPR58[31] , 
        \B_DOUT_TEMPR59[31] , \B_DOUT_TEMPR60[31] , 
        \B_DOUT_TEMPR61[31] , \B_DOUT_TEMPR62[31] , 
        \B_DOUT_TEMPR63[31] , \B_DOUT_TEMPR64[31] , 
        \B_DOUT_TEMPR65[31] , \B_DOUT_TEMPR66[31] , 
        \B_DOUT_TEMPR67[31] , \B_DOUT_TEMPR68[31] , 
        \B_DOUT_TEMPR69[31] , \B_DOUT_TEMPR70[31] , 
        \B_DOUT_TEMPR71[31] , \B_DOUT_TEMPR72[31] , 
        \B_DOUT_TEMPR73[31] , \B_DOUT_TEMPR74[31] , 
        \B_DOUT_TEMPR75[31] , \B_DOUT_TEMPR76[31] , 
        \B_DOUT_TEMPR77[31] , \B_DOUT_TEMPR78[31] , 
        \B_DOUT_TEMPR79[31] , \B_DOUT_TEMPR80[31] , 
        \B_DOUT_TEMPR81[31] , \B_DOUT_TEMPR82[31] , 
        \B_DOUT_TEMPR83[31] , \B_DOUT_TEMPR84[31] , 
        \B_DOUT_TEMPR85[31] , \B_DOUT_TEMPR86[31] , 
        \B_DOUT_TEMPR87[31] , \B_DOUT_TEMPR88[31] , 
        \B_DOUT_TEMPR89[31] , \B_DOUT_TEMPR90[31] , 
        \B_DOUT_TEMPR91[31] , \B_DOUT_TEMPR92[31] , 
        \B_DOUT_TEMPR93[31] , \B_DOUT_TEMPR94[31] , 
        \B_DOUT_TEMPR95[31] , \B_DOUT_TEMPR96[31] , 
        \B_DOUT_TEMPR97[31] , \B_DOUT_TEMPR98[31] , 
        \B_DOUT_TEMPR99[31] , \B_DOUT_TEMPR100[31] , 
        \B_DOUT_TEMPR101[31] , \B_DOUT_TEMPR102[31] , 
        \B_DOUT_TEMPR103[31] , \B_DOUT_TEMPR104[31] , 
        \B_DOUT_TEMPR105[31] , \B_DOUT_TEMPR106[31] , 
        \B_DOUT_TEMPR107[31] , \B_DOUT_TEMPR108[31] , 
        \B_DOUT_TEMPR109[31] , \B_DOUT_TEMPR110[31] , 
        \B_DOUT_TEMPR111[31] , \B_DOUT_TEMPR112[31] , 
        \B_DOUT_TEMPR113[31] , \B_DOUT_TEMPR114[31] , 
        \B_DOUT_TEMPR115[31] , \B_DOUT_TEMPR116[31] , 
        \B_DOUT_TEMPR117[31] , \B_DOUT_TEMPR118[31] , 
        \B_DOUT_TEMPR0[32] , \B_DOUT_TEMPR1[32] , \B_DOUT_TEMPR2[32] , 
        \B_DOUT_TEMPR3[32] , \B_DOUT_TEMPR4[32] , \B_DOUT_TEMPR5[32] , 
        \B_DOUT_TEMPR6[32] , \B_DOUT_TEMPR7[32] , \B_DOUT_TEMPR8[32] , 
        \B_DOUT_TEMPR9[32] , \B_DOUT_TEMPR10[32] , 
        \B_DOUT_TEMPR11[32] , \B_DOUT_TEMPR12[32] , 
        \B_DOUT_TEMPR13[32] , \B_DOUT_TEMPR14[32] , 
        \B_DOUT_TEMPR15[32] , \B_DOUT_TEMPR16[32] , 
        \B_DOUT_TEMPR17[32] , \B_DOUT_TEMPR18[32] , 
        \B_DOUT_TEMPR19[32] , \B_DOUT_TEMPR20[32] , 
        \B_DOUT_TEMPR21[32] , \B_DOUT_TEMPR22[32] , 
        \B_DOUT_TEMPR23[32] , \B_DOUT_TEMPR24[32] , 
        \B_DOUT_TEMPR25[32] , \B_DOUT_TEMPR26[32] , 
        \B_DOUT_TEMPR27[32] , \B_DOUT_TEMPR28[32] , 
        \B_DOUT_TEMPR29[32] , \B_DOUT_TEMPR30[32] , 
        \B_DOUT_TEMPR31[32] , \B_DOUT_TEMPR32[32] , 
        \B_DOUT_TEMPR33[32] , \B_DOUT_TEMPR34[32] , 
        \B_DOUT_TEMPR35[32] , \B_DOUT_TEMPR36[32] , 
        \B_DOUT_TEMPR37[32] , \B_DOUT_TEMPR38[32] , 
        \B_DOUT_TEMPR39[32] , \B_DOUT_TEMPR40[32] , 
        \B_DOUT_TEMPR41[32] , \B_DOUT_TEMPR42[32] , 
        \B_DOUT_TEMPR43[32] , \B_DOUT_TEMPR44[32] , 
        \B_DOUT_TEMPR45[32] , \B_DOUT_TEMPR46[32] , 
        \B_DOUT_TEMPR47[32] , \B_DOUT_TEMPR48[32] , 
        \B_DOUT_TEMPR49[32] , \B_DOUT_TEMPR50[32] , 
        \B_DOUT_TEMPR51[32] , \B_DOUT_TEMPR52[32] , 
        \B_DOUT_TEMPR53[32] , \B_DOUT_TEMPR54[32] , 
        \B_DOUT_TEMPR55[32] , \B_DOUT_TEMPR56[32] , 
        \B_DOUT_TEMPR57[32] , \B_DOUT_TEMPR58[32] , 
        \B_DOUT_TEMPR59[32] , \B_DOUT_TEMPR60[32] , 
        \B_DOUT_TEMPR61[32] , \B_DOUT_TEMPR62[32] , 
        \B_DOUT_TEMPR63[32] , \B_DOUT_TEMPR64[32] , 
        \B_DOUT_TEMPR65[32] , \B_DOUT_TEMPR66[32] , 
        \B_DOUT_TEMPR67[32] , \B_DOUT_TEMPR68[32] , 
        \B_DOUT_TEMPR69[32] , \B_DOUT_TEMPR70[32] , 
        \B_DOUT_TEMPR71[32] , \B_DOUT_TEMPR72[32] , 
        \B_DOUT_TEMPR73[32] , \B_DOUT_TEMPR74[32] , 
        \B_DOUT_TEMPR75[32] , \B_DOUT_TEMPR76[32] , 
        \B_DOUT_TEMPR77[32] , \B_DOUT_TEMPR78[32] , 
        \B_DOUT_TEMPR79[32] , \B_DOUT_TEMPR80[32] , 
        \B_DOUT_TEMPR81[32] , \B_DOUT_TEMPR82[32] , 
        \B_DOUT_TEMPR83[32] , \B_DOUT_TEMPR84[32] , 
        \B_DOUT_TEMPR85[32] , \B_DOUT_TEMPR86[32] , 
        \B_DOUT_TEMPR87[32] , \B_DOUT_TEMPR88[32] , 
        \B_DOUT_TEMPR89[32] , \B_DOUT_TEMPR90[32] , 
        \B_DOUT_TEMPR91[32] , \B_DOUT_TEMPR92[32] , 
        \B_DOUT_TEMPR93[32] , \B_DOUT_TEMPR94[32] , 
        \B_DOUT_TEMPR95[32] , \B_DOUT_TEMPR96[32] , 
        \B_DOUT_TEMPR97[32] , \B_DOUT_TEMPR98[32] , 
        \B_DOUT_TEMPR99[32] , \B_DOUT_TEMPR100[32] , 
        \B_DOUT_TEMPR101[32] , \B_DOUT_TEMPR102[32] , 
        \B_DOUT_TEMPR103[32] , \B_DOUT_TEMPR104[32] , 
        \B_DOUT_TEMPR105[32] , \B_DOUT_TEMPR106[32] , 
        \B_DOUT_TEMPR107[32] , \B_DOUT_TEMPR108[32] , 
        \B_DOUT_TEMPR109[32] , \B_DOUT_TEMPR110[32] , 
        \B_DOUT_TEMPR111[32] , \B_DOUT_TEMPR112[32] , 
        \B_DOUT_TEMPR113[32] , \B_DOUT_TEMPR114[32] , 
        \B_DOUT_TEMPR115[32] , \B_DOUT_TEMPR116[32] , 
        \B_DOUT_TEMPR117[32] , \B_DOUT_TEMPR118[32] , 
        \B_DOUT_TEMPR0[33] , \B_DOUT_TEMPR1[33] , \B_DOUT_TEMPR2[33] , 
        \B_DOUT_TEMPR3[33] , \B_DOUT_TEMPR4[33] , \B_DOUT_TEMPR5[33] , 
        \B_DOUT_TEMPR6[33] , \B_DOUT_TEMPR7[33] , \B_DOUT_TEMPR8[33] , 
        \B_DOUT_TEMPR9[33] , \B_DOUT_TEMPR10[33] , 
        \B_DOUT_TEMPR11[33] , \B_DOUT_TEMPR12[33] , 
        \B_DOUT_TEMPR13[33] , \B_DOUT_TEMPR14[33] , 
        \B_DOUT_TEMPR15[33] , \B_DOUT_TEMPR16[33] , 
        \B_DOUT_TEMPR17[33] , \B_DOUT_TEMPR18[33] , 
        \B_DOUT_TEMPR19[33] , \B_DOUT_TEMPR20[33] , 
        \B_DOUT_TEMPR21[33] , \B_DOUT_TEMPR22[33] , 
        \B_DOUT_TEMPR23[33] , \B_DOUT_TEMPR24[33] , 
        \B_DOUT_TEMPR25[33] , \B_DOUT_TEMPR26[33] , 
        \B_DOUT_TEMPR27[33] , \B_DOUT_TEMPR28[33] , 
        \B_DOUT_TEMPR29[33] , \B_DOUT_TEMPR30[33] , 
        \B_DOUT_TEMPR31[33] , \B_DOUT_TEMPR32[33] , 
        \B_DOUT_TEMPR33[33] , \B_DOUT_TEMPR34[33] , 
        \B_DOUT_TEMPR35[33] , \B_DOUT_TEMPR36[33] , 
        \B_DOUT_TEMPR37[33] , \B_DOUT_TEMPR38[33] , 
        \B_DOUT_TEMPR39[33] , \B_DOUT_TEMPR40[33] , 
        \B_DOUT_TEMPR41[33] , \B_DOUT_TEMPR42[33] , 
        \B_DOUT_TEMPR43[33] , \B_DOUT_TEMPR44[33] , 
        \B_DOUT_TEMPR45[33] , \B_DOUT_TEMPR46[33] , 
        \B_DOUT_TEMPR47[33] , \B_DOUT_TEMPR48[33] , 
        \B_DOUT_TEMPR49[33] , \B_DOUT_TEMPR50[33] , 
        \B_DOUT_TEMPR51[33] , \B_DOUT_TEMPR52[33] , 
        \B_DOUT_TEMPR53[33] , \B_DOUT_TEMPR54[33] , 
        \B_DOUT_TEMPR55[33] , \B_DOUT_TEMPR56[33] , 
        \B_DOUT_TEMPR57[33] , \B_DOUT_TEMPR58[33] , 
        \B_DOUT_TEMPR59[33] , \B_DOUT_TEMPR60[33] , 
        \B_DOUT_TEMPR61[33] , \B_DOUT_TEMPR62[33] , 
        \B_DOUT_TEMPR63[33] , \B_DOUT_TEMPR64[33] , 
        \B_DOUT_TEMPR65[33] , \B_DOUT_TEMPR66[33] , 
        \B_DOUT_TEMPR67[33] , \B_DOUT_TEMPR68[33] , 
        \B_DOUT_TEMPR69[33] , \B_DOUT_TEMPR70[33] , 
        \B_DOUT_TEMPR71[33] , \B_DOUT_TEMPR72[33] , 
        \B_DOUT_TEMPR73[33] , \B_DOUT_TEMPR74[33] , 
        \B_DOUT_TEMPR75[33] , \B_DOUT_TEMPR76[33] , 
        \B_DOUT_TEMPR77[33] , \B_DOUT_TEMPR78[33] , 
        \B_DOUT_TEMPR79[33] , \B_DOUT_TEMPR80[33] , 
        \B_DOUT_TEMPR81[33] , \B_DOUT_TEMPR82[33] , 
        \B_DOUT_TEMPR83[33] , \B_DOUT_TEMPR84[33] , 
        \B_DOUT_TEMPR85[33] , \B_DOUT_TEMPR86[33] , 
        \B_DOUT_TEMPR87[33] , \B_DOUT_TEMPR88[33] , 
        \B_DOUT_TEMPR89[33] , \B_DOUT_TEMPR90[33] , 
        \B_DOUT_TEMPR91[33] , \B_DOUT_TEMPR92[33] , 
        \B_DOUT_TEMPR93[33] , \B_DOUT_TEMPR94[33] , 
        \B_DOUT_TEMPR95[33] , \B_DOUT_TEMPR96[33] , 
        \B_DOUT_TEMPR97[33] , \B_DOUT_TEMPR98[33] , 
        \B_DOUT_TEMPR99[33] , \B_DOUT_TEMPR100[33] , 
        \B_DOUT_TEMPR101[33] , \B_DOUT_TEMPR102[33] , 
        \B_DOUT_TEMPR103[33] , \B_DOUT_TEMPR104[33] , 
        \B_DOUT_TEMPR105[33] , \B_DOUT_TEMPR106[33] , 
        \B_DOUT_TEMPR107[33] , \B_DOUT_TEMPR108[33] , 
        \B_DOUT_TEMPR109[33] , \B_DOUT_TEMPR110[33] , 
        \B_DOUT_TEMPR111[33] , \B_DOUT_TEMPR112[33] , 
        \B_DOUT_TEMPR113[33] , \B_DOUT_TEMPR114[33] , 
        \B_DOUT_TEMPR115[33] , \B_DOUT_TEMPR116[33] , 
        \B_DOUT_TEMPR117[33] , \B_DOUT_TEMPR118[33] , 
        \B_DOUT_TEMPR0[34] , \B_DOUT_TEMPR1[34] , \B_DOUT_TEMPR2[34] , 
        \B_DOUT_TEMPR3[34] , \B_DOUT_TEMPR4[34] , \B_DOUT_TEMPR5[34] , 
        \B_DOUT_TEMPR6[34] , \B_DOUT_TEMPR7[34] , \B_DOUT_TEMPR8[34] , 
        \B_DOUT_TEMPR9[34] , \B_DOUT_TEMPR10[34] , 
        \B_DOUT_TEMPR11[34] , \B_DOUT_TEMPR12[34] , 
        \B_DOUT_TEMPR13[34] , \B_DOUT_TEMPR14[34] , 
        \B_DOUT_TEMPR15[34] , \B_DOUT_TEMPR16[34] , 
        \B_DOUT_TEMPR17[34] , \B_DOUT_TEMPR18[34] , 
        \B_DOUT_TEMPR19[34] , \B_DOUT_TEMPR20[34] , 
        \B_DOUT_TEMPR21[34] , \B_DOUT_TEMPR22[34] , 
        \B_DOUT_TEMPR23[34] , \B_DOUT_TEMPR24[34] , 
        \B_DOUT_TEMPR25[34] , \B_DOUT_TEMPR26[34] , 
        \B_DOUT_TEMPR27[34] , \B_DOUT_TEMPR28[34] , 
        \B_DOUT_TEMPR29[34] , \B_DOUT_TEMPR30[34] , 
        \B_DOUT_TEMPR31[34] , \B_DOUT_TEMPR32[34] , 
        \B_DOUT_TEMPR33[34] , \B_DOUT_TEMPR34[34] , 
        \B_DOUT_TEMPR35[34] , \B_DOUT_TEMPR36[34] , 
        \B_DOUT_TEMPR37[34] , \B_DOUT_TEMPR38[34] , 
        \B_DOUT_TEMPR39[34] , \B_DOUT_TEMPR40[34] , 
        \B_DOUT_TEMPR41[34] , \B_DOUT_TEMPR42[34] , 
        \B_DOUT_TEMPR43[34] , \B_DOUT_TEMPR44[34] , 
        \B_DOUT_TEMPR45[34] , \B_DOUT_TEMPR46[34] , 
        \B_DOUT_TEMPR47[34] , \B_DOUT_TEMPR48[34] , 
        \B_DOUT_TEMPR49[34] , \B_DOUT_TEMPR50[34] , 
        \B_DOUT_TEMPR51[34] , \B_DOUT_TEMPR52[34] , 
        \B_DOUT_TEMPR53[34] , \B_DOUT_TEMPR54[34] , 
        \B_DOUT_TEMPR55[34] , \B_DOUT_TEMPR56[34] , 
        \B_DOUT_TEMPR57[34] , \B_DOUT_TEMPR58[34] , 
        \B_DOUT_TEMPR59[34] , \B_DOUT_TEMPR60[34] , 
        \B_DOUT_TEMPR61[34] , \B_DOUT_TEMPR62[34] , 
        \B_DOUT_TEMPR63[34] , \B_DOUT_TEMPR64[34] , 
        \B_DOUT_TEMPR65[34] , \B_DOUT_TEMPR66[34] , 
        \B_DOUT_TEMPR67[34] , \B_DOUT_TEMPR68[34] , 
        \B_DOUT_TEMPR69[34] , \B_DOUT_TEMPR70[34] , 
        \B_DOUT_TEMPR71[34] , \B_DOUT_TEMPR72[34] , 
        \B_DOUT_TEMPR73[34] , \B_DOUT_TEMPR74[34] , 
        \B_DOUT_TEMPR75[34] , \B_DOUT_TEMPR76[34] , 
        \B_DOUT_TEMPR77[34] , \B_DOUT_TEMPR78[34] , 
        \B_DOUT_TEMPR79[34] , \B_DOUT_TEMPR80[34] , 
        \B_DOUT_TEMPR81[34] , \B_DOUT_TEMPR82[34] , 
        \B_DOUT_TEMPR83[34] , \B_DOUT_TEMPR84[34] , 
        \B_DOUT_TEMPR85[34] , \B_DOUT_TEMPR86[34] , 
        \B_DOUT_TEMPR87[34] , \B_DOUT_TEMPR88[34] , 
        \B_DOUT_TEMPR89[34] , \B_DOUT_TEMPR90[34] , 
        \B_DOUT_TEMPR91[34] , \B_DOUT_TEMPR92[34] , 
        \B_DOUT_TEMPR93[34] , \B_DOUT_TEMPR94[34] , 
        \B_DOUT_TEMPR95[34] , \B_DOUT_TEMPR96[34] , 
        \B_DOUT_TEMPR97[34] , \B_DOUT_TEMPR98[34] , 
        \B_DOUT_TEMPR99[34] , \B_DOUT_TEMPR100[34] , 
        \B_DOUT_TEMPR101[34] , \B_DOUT_TEMPR102[34] , 
        \B_DOUT_TEMPR103[34] , \B_DOUT_TEMPR104[34] , 
        \B_DOUT_TEMPR105[34] , \B_DOUT_TEMPR106[34] , 
        \B_DOUT_TEMPR107[34] , \B_DOUT_TEMPR108[34] , 
        \B_DOUT_TEMPR109[34] , \B_DOUT_TEMPR110[34] , 
        \B_DOUT_TEMPR111[34] , \B_DOUT_TEMPR112[34] , 
        \B_DOUT_TEMPR113[34] , \B_DOUT_TEMPR114[34] , 
        \B_DOUT_TEMPR115[34] , \B_DOUT_TEMPR116[34] , 
        \B_DOUT_TEMPR117[34] , \B_DOUT_TEMPR118[34] , 
        \B_DOUT_TEMPR0[35] , \B_DOUT_TEMPR1[35] , \B_DOUT_TEMPR2[35] , 
        \B_DOUT_TEMPR3[35] , \B_DOUT_TEMPR4[35] , \B_DOUT_TEMPR5[35] , 
        \B_DOUT_TEMPR6[35] , \B_DOUT_TEMPR7[35] , \B_DOUT_TEMPR8[35] , 
        \B_DOUT_TEMPR9[35] , \B_DOUT_TEMPR10[35] , 
        \B_DOUT_TEMPR11[35] , \B_DOUT_TEMPR12[35] , 
        \B_DOUT_TEMPR13[35] , \B_DOUT_TEMPR14[35] , 
        \B_DOUT_TEMPR15[35] , \B_DOUT_TEMPR16[35] , 
        \B_DOUT_TEMPR17[35] , \B_DOUT_TEMPR18[35] , 
        \B_DOUT_TEMPR19[35] , \B_DOUT_TEMPR20[35] , 
        \B_DOUT_TEMPR21[35] , \B_DOUT_TEMPR22[35] , 
        \B_DOUT_TEMPR23[35] , \B_DOUT_TEMPR24[35] , 
        \B_DOUT_TEMPR25[35] , \B_DOUT_TEMPR26[35] , 
        \B_DOUT_TEMPR27[35] , \B_DOUT_TEMPR28[35] , 
        \B_DOUT_TEMPR29[35] , \B_DOUT_TEMPR30[35] , 
        \B_DOUT_TEMPR31[35] , \B_DOUT_TEMPR32[35] , 
        \B_DOUT_TEMPR33[35] , \B_DOUT_TEMPR34[35] , 
        \B_DOUT_TEMPR35[35] , \B_DOUT_TEMPR36[35] , 
        \B_DOUT_TEMPR37[35] , \B_DOUT_TEMPR38[35] , 
        \B_DOUT_TEMPR39[35] , \B_DOUT_TEMPR40[35] , 
        \B_DOUT_TEMPR41[35] , \B_DOUT_TEMPR42[35] , 
        \B_DOUT_TEMPR43[35] , \B_DOUT_TEMPR44[35] , 
        \B_DOUT_TEMPR45[35] , \B_DOUT_TEMPR46[35] , 
        \B_DOUT_TEMPR47[35] , \B_DOUT_TEMPR48[35] , 
        \B_DOUT_TEMPR49[35] , \B_DOUT_TEMPR50[35] , 
        \B_DOUT_TEMPR51[35] , \B_DOUT_TEMPR52[35] , 
        \B_DOUT_TEMPR53[35] , \B_DOUT_TEMPR54[35] , 
        \B_DOUT_TEMPR55[35] , \B_DOUT_TEMPR56[35] , 
        \B_DOUT_TEMPR57[35] , \B_DOUT_TEMPR58[35] , 
        \B_DOUT_TEMPR59[35] , \B_DOUT_TEMPR60[35] , 
        \B_DOUT_TEMPR61[35] , \B_DOUT_TEMPR62[35] , 
        \B_DOUT_TEMPR63[35] , \B_DOUT_TEMPR64[35] , 
        \B_DOUT_TEMPR65[35] , \B_DOUT_TEMPR66[35] , 
        \B_DOUT_TEMPR67[35] , \B_DOUT_TEMPR68[35] , 
        \B_DOUT_TEMPR69[35] , \B_DOUT_TEMPR70[35] , 
        \B_DOUT_TEMPR71[35] , \B_DOUT_TEMPR72[35] , 
        \B_DOUT_TEMPR73[35] , \B_DOUT_TEMPR74[35] , 
        \B_DOUT_TEMPR75[35] , \B_DOUT_TEMPR76[35] , 
        \B_DOUT_TEMPR77[35] , \B_DOUT_TEMPR78[35] , 
        \B_DOUT_TEMPR79[35] , \B_DOUT_TEMPR80[35] , 
        \B_DOUT_TEMPR81[35] , \B_DOUT_TEMPR82[35] , 
        \B_DOUT_TEMPR83[35] , \B_DOUT_TEMPR84[35] , 
        \B_DOUT_TEMPR85[35] , \B_DOUT_TEMPR86[35] , 
        \B_DOUT_TEMPR87[35] , \B_DOUT_TEMPR88[35] , 
        \B_DOUT_TEMPR89[35] , \B_DOUT_TEMPR90[35] , 
        \B_DOUT_TEMPR91[35] , \B_DOUT_TEMPR92[35] , 
        \B_DOUT_TEMPR93[35] , \B_DOUT_TEMPR94[35] , 
        \B_DOUT_TEMPR95[35] , \B_DOUT_TEMPR96[35] , 
        \B_DOUT_TEMPR97[35] , \B_DOUT_TEMPR98[35] , 
        \B_DOUT_TEMPR99[35] , \B_DOUT_TEMPR100[35] , 
        \B_DOUT_TEMPR101[35] , \B_DOUT_TEMPR102[35] , 
        \B_DOUT_TEMPR103[35] , \B_DOUT_TEMPR104[35] , 
        \B_DOUT_TEMPR105[35] , \B_DOUT_TEMPR106[35] , 
        \B_DOUT_TEMPR107[35] , \B_DOUT_TEMPR108[35] , 
        \B_DOUT_TEMPR109[35] , \B_DOUT_TEMPR110[35] , 
        \B_DOUT_TEMPR111[35] , \B_DOUT_TEMPR112[35] , 
        \B_DOUT_TEMPR113[35] , \B_DOUT_TEMPR114[35] , 
        \B_DOUT_TEMPR115[35] , \B_DOUT_TEMPR116[35] , 
        \B_DOUT_TEMPR117[35] , \B_DOUT_TEMPR118[35] , 
        \B_DOUT_TEMPR0[36] , \B_DOUT_TEMPR1[36] , \B_DOUT_TEMPR2[36] , 
        \B_DOUT_TEMPR3[36] , \B_DOUT_TEMPR4[36] , \B_DOUT_TEMPR5[36] , 
        \B_DOUT_TEMPR6[36] , \B_DOUT_TEMPR7[36] , \B_DOUT_TEMPR8[36] , 
        \B_DOUT_TEMPR9[36] , \B_DOUT_TEMPR10[36] , 
        \B_DOUT_TEMPR11[36] , \B_DOUT_TEMPR12[36] , 
        \B_DOUT_TEMPR13[36] , \B_DOUT_TEMPR14[36] , 
        \B_DOUT_TEMPR15[36] , \B_DOUT_TEMPR16[36] , 
        \B_DOUT_TEMPR17[36] , \B_DOUT_TEMPR18[36] , 
        \B_DOUT_TEMPR19[36] , \B_DOUT_TEMPR20[36] , 
        \B_DOUT_TEMPR21[36] , \B_DOUT_TEMPR22[36] , 
        \B_DOUT_TEMPR23[36] , \B_DOUT_TEMPR24[36] , 
        \B_DOUT_TEMPR25[36] , \B_DOUT_TEMPR26[36] , 
        \B_DOUT_TEMPR27[36] , \B_DOUT_TEMPR28[36] , 
        \B_DOUT_TEMPR29[36] , \B_DOUT_TEMPR30[36] , 
        \B_DOUT_TEMPR31[36] , \B_DOUT_TEMPR32[36] , 
        \B_DOUT_TEMPR33[36] , \B_DOUT_TEMPR34[36] , 
        \B_DOUT_TEMPR35[36] , \B_DOUT_TEMPR36[36] , 
        \B_DOUT_TEMPR37[36] , \B_DOUT_TEMPR38[36] , 
        \B_DOUT_TEMPR39[36] , \B_DOUT_TEMPR40[36] , 
        \B_DOUT_TEMPR41[36] , \B_DOUT_TEMPR42[36] , 
        \B_DOUT_TEMPR43[36] , \B_DOUT_TEMPR44[36] , 
        \B_DOUT_TEMPR45[36] , \B_DOUT_TEMPR46[36] , 
        \B_DOUT_TEMPR47[36] , \B_DOUT_TEMPR48[36] , 
        \B_DOUT_TEMPR49[36] , \B_DOUT_TEMPR50[36] , 
        \B_DOUT_TEMPR51[36] , \B_DOUT_TEMPR52[36] , 
        \B_DOUT_TEMPR53[36] , \B_DOUT_TEMPR54[36] , 
        \B_DOUT_TEMPR55[36] , \B_DOUT_TEMPR56[36] , 
        \B_DOUT_TEMPR57[36] , \B_DOUT_TEMPR58[36] , 
        \B_DOUT_TEMPR59[36] , \B_DOUT_TEMPR60[36] , 
        \B_DOUT_TEMPR61[36] , \B_DOUT_TEMPR62[36] , 
        \B_DOUT_TEMPR63[36] , \B_DOUT_TEMPR64[36] , 
        \B_DOUT_TEMPR65[36] , \B_DOUT_TEMPR66[36] , 
        \B_DOUT_TEMPR67[36] , \B_DOUT_TEMPR68[36] , 
        \B_DOUT_TEMPR69[36] , \B_DOUT_TEMPR70[36] , 
        \B_DOUT_TEMPR71[36] , \B_DOUT_TEMPR72[36] , 
        \B_DOUT_TEMPR73[36] , \B_DOUT_TEMPR74[36] , 
        \B_DOUT_TEMPR75[36] , \B_DOUT_TEMPR76[36] , 
        \B_DOUT_TEMPR77[36] , \B_DOUT_TEMPR78[36] , 
        \B_DOUT_TEMPR79[36] , \B_DOUT_TEMPR80[36] , 
        \B_DOUT_TEMPR81[36] , \B_DOUT_TEMPR82[36] , 
        \B_DOUT_TEMPR83[36] , \B_DOUT_TEMPR84[36] , 
        \B_DOUT_TEMPR85[36] , \B_DOUT_TEMPR86[36] , 
        \B_DOUT_TEMPR87[36] , \B_DOUT_TEMPR88[36] , 
        \B_DOUT_TEMPR89[36] , \B_DOUT_TEMPR90[36] , 
        \B_DOUT_TEMPR91[36] , \B_DOUT_TEMPR92[36] , 
        \B_DOUT_TEMPR93[36] , \B_DOUT_TEMPR94[36] , 
        \B_DOUT_TEMPR95[36] , \B_DOUT_TEMPR96[36] , 
        \B_DOUT_TEMPR97[36] , \B_DOUT_TEMPR98[36] , 
        \B_DOUT_TEMPR99[36] , \B_DOUT_TEMPR100[36] , 
        \B_DOUT_TEMPR101[36] , \B_DOUT_TEMPR102[36] , 
        \B_DOUT_TEMPR103[36] , \B_DOUT_TEMPR104[36] , 
        \B_DOUT_TEMPR105[36] , \B_DOUT_TEMPR106[36] , 
        \B_DOUT_TEMPR107[36] , \B_DOUT_TEMPR108[36] , 
        \B_DOUT_TEMPR109[36] , \B_DOUT_TEMPR110[36] , 
        \B_DOUT_TEMPR111[36] , \B_DOUT_TEMPR112[36] , 
        \B_DOUT_TEMPR113[36] , \B_DOUT_TEMPR114[36] , 
        \B_DOUT_TEMPR115[36] , \B_DOUT_TEMPR116[36] , 
        \B_DOUT_TEMPR117[36] , \B_DOUT_TEMPR118[36] , 
        \B_DOUT_TEMPR0[37] , \B_DOUT_TEMPR1[37] , \B_DOUT_TEMPR2[37] , 
        \B_DOUT_TEMPR3[37] , \B_DOUT_TEMPR4[37] , \B_DOUT_TEMPR5[37] , 
        \B_DOUT_TEMPR6[37] , \B_DOUT_TEMPR7[37] , \B_DOUT_TEMPR8[37] , 
        \B_DOUT_TEMPR9[37] , \B_DOUT_TEMPR10[37] , 
        \B_DOUT_TEMPR11[37] , \B_DOUT_TEMPR12[37] , 
        \B_DOUT_TEMPR13[37] , \B_DOUT_TEMPR14[37] , 
        \B_DOUT_TEMPR15[37] , \B_DOUT_TEMPR16[37] , 
        \B_DOUT_TEMPR17[37] , \B_DOUT_TEMPR18[37] , 
        \B_DOUT_TEMPR19[37] , \B_DOUT_TEMPR20[37] , 
        \B_DOUT_TEMPR21[37] , \B_DOUT_TEMPR22[37] , 
        \B_DOUT_TEMPR23[37] , \B_DOUT_TEMPR24[37] , 
        \B_DOUT_TEMPR25[37] , \B_DOUT_TEMPR26[37] , 
        \B_DOUT_TEMPR27[37] , \B_DOUT_TEMPR28[37] , 
        \B_DOUT_TEMPR29[37] , \B_DOUT_TEMPR30[37] , 
        \B_DOUT_TEMPR31[37] , \B_DOUT_TEMPR32[37] , 
        \B_DOUT_TEMPR33[37] , \B_DOUT_TEMPR34[37] , 
        \B_DOUT_TEMPR35[37] , \B_DOUT_TEMPR36[37] , 
        \B_DOUT_TEMPR37[37] , \B_DOUT_TEMPR38[37] , 
        \B_DOUT_TEMPR39[37] , \B_DOUT_TEMPR40[37] , 
        \B_DOUT_TEMPR41[37] , \B_DOUT_TEMPR42[37] , 
        \B_DOUT_TEMPR43[37] , \B_DOUT_TEMPR44[37] , 
        \B_DOUT_TEMPR45[37] , \B_DOUT_TEMPR46[37] , 
        \B_DOUT_TEMPR47[37] , \B_DOUT_TEMPR48[37] , 
        \B_DOUT_TEMPR49[37] , \B_DOUT_TEMPR50[37] , 
        \B_DOUT_TEMPR51[37] , \B_DOUT_TEMPR52[37] , 
        \B_DOUT_TEMPR53[37] , \B_DOUT_TEMPR54[37] , 
        \B_DOUT_TEMPR55[37] , \B_DOUT_TEMPR56[37] , 
        \B_DOUT_TEMPR57[37] , \B_DOUT_TEMPR58[37] , 
        \B_DOUT_TEMPR59[37] , \B_DOUT_TEMPR60[37] , 
        \B_DOUT_TEMPR61[37] , \B_DOUT_TEMPR62[37] , 
        \B_DOUT_TEMPR63[37] , \B_DOUT_TEMPR64[37] , 
        \B_DOUT_TEMPR65[37] , \B_DOUT_TEMPR66[37] , 
        \B_DOUT_TEMPR67[37] , \B_DOUT_TEMPR68[37] , 
        \B_DOUT_TEMPR69[37] , \B_DOUT_TEMPR70[37] , 
        \B_DOUT_TEMPR71[37] , \B_DOUT_TEMPR72[37] , 
        \B_DOUT_TEMPR73[37] , \B_DOUT_TEMPR74[37] , 
        \B_DOUT_TEMPR75[37] , \B_DOUT_TEMPR76[37] , 
        \B_DOUT_TEMPR77[37] , \B_DOUT_TEMPR78[37] , 
        \B_DOUT_TEMPR79[37] , \B_DOUT_TEMPR80[37] , 
        \B_DOUT_TEMPR81[37] , \B_DOUT_TEMPR82[37] , 
        \B_DOUT_TEMPR83[37] , \B_DOUT_TEMPR84[37] , 
        \B_DOUT_TEMPR85[37] , \B_DOUT_TEMPR86[37] , 
        \B_DOUT_TEMPR87[37] , \B_DOUT_TEMPR88[37] , 
        \B_DOUT_TEMPR89[37] , \B_DOUT_TEMPR90[37] , 
        \B_DOUT_TEMPR91[37] , \B_DOUT_TEMPR92[37] , 
        \B_DOUT_TEMPR93[37] , \B_DOUT_TEMPR94[37] , 
        \B_DOUT_TEMPR95[37] , \B_DOUT_TEMPR96[37] , 
        \B_DOUT_TEMPR97[37] , \B_DOUT_TEMPR98[37] , 
        \B_DOUT_TEMPR99[37] , \B_DOUT_TEMPR100[37] , 
        \B_DOUT_TEMPR101[37] , \B_DOUT_TEMPR102[37] , 
        \B_DOUT_TEMPR103[37] , \B_DOUT_TEMPR104[37] , 
        \B_DOUT_TEMPR105[37] , \B_DOUT_TEMPR106[37] , 
        \B_DOUT_TEMPR107[37] , \B_DOUT_TEMPR108[37] , 
        \B_DOUT_TEMPR109[37] , \B_DOUT_TEMPR110[37] , 
        \B_DOUT_TEMPR111[37] , \B_DOUT_TEMPR112[37] , 
        \B_DOUT_TEMPR113[37] , \B_DOUT_TEMPR114[37] , 
        \B_DOUT_TEMPR115[37] , \B_DOUT_TEMPR116[37] , 
        \B_DOUT_TEMPR117[37] , \B_DOUT_TEMPR118[37] , 
        \B_DOUT_TEMPR0[38] , \B_DOUT_TEMPR1[38] , \B_DOUT_TEMPR2[38] , 
        \B_DOUT_TEMPR3[38] , \B_DOUT_TEMPR4[38] , \B_DOUT_TEMPR5[38] , 
        \B_DOUT_TEMPR6[38] , \B_DOUT_TEMPR7[38] , \B_DOUT_TEMPR8[38] , 
        \B_DOUT_TEMPR9[38] , \B_DOUT_TEMPR10[38] , 
        \B_DOUT_TEMPR11[38] , \B_DOUT_TEMPR12[38] , 
        \B_DOUT_TEMPR13[38] , \B_DOUT_TEMPR14[38] , 
        \B_DOUT_TEMPR15[38] , \B_DOUT_TEMPR16[38] , 
        \B_DOUT_TEMPR17[38] , \B_DOUT_TEMPR18[38] , 
        \B_DOUT_TEMPR19[38] , \B_DOUT_TEMPR20[38] , 
        \B_DOUT_TEMPR21[38] , \B_DOUT_TEMPR22[38] , 
        \B_DOUT_TEMPR23[38] , \B_DOUT_TEMPR24[38] , 
        \B_DOUT_TEMPR25[38] , \B_DOUT_TEMPR26[38] , 
        \B_DOUT_TEMPR27[38] , \B_DOUT_TEMPR28[38] , 
        \B_DOUT_TEMPR29[38] , \B_DOUT_TEMPR30[38] , 
        \B_DOUT_TEMPR31[38] , \B_DOUT_TEMPR32[38] , 
        \B_DOUT_TEMPR33[38] , \B_DOUT_TEMPR34[38] , 
        \B_DOUT_TEMPR35[38] , \B_DOUT_TEMPR36[38] , 
        \B_DOUT_TEMPR37[38] , \B_DOUT_TEMPR38[38] , 
        \B_DOUT_TEMPR39[38] , \B_DOUT_TEMPR40[38] , 
        \B_DOUT_TEMPR41[38] , \B_DOUT_TEMPR42[38] , 
        \B_DOUT_TEMPR43[38] , \B_DOUT_TEMPR44[38] , 
        \B_DOUT_TEMPR45[38] , \B_DOUT_TEMPR46[38] , 
        \B_DOUT_TEMPR47[38] , \B_DOUT_TEMPR48[38] , 
        \B_DOUT_TEMPR49[38] , \B_DOUT_TEMPR50[38] , 
        \B_DOUT_TEMPR51[38] , \B_DOUT_TEMPR52[38] , 
        \B_DOUT_TEMPR53[38] , \B_DOUT_TEMPR54[38] , 
        \B_DOUT_TEMPR55[38] , \B_DOUT_TEMPR56[38] , 
        \B_DOUT_TEMPR57[38] , \B_DOUT_TEMPR58[38] , 
        \B_DOUT_TEMPR59[38] , \B_DOUT_TEMPR60[38] , 
        \B_DOUT_TEMPR61[38] , \B_DOUT_TEMPR62[38] , 
        \B_DOUT_TEMPR63[38] , \B_DOUT_TEMPR64[38] , 
        \B_DOUT_TEMPR65[38] , \B_DOUT_TEMPR66[38] , 
        \B_DOUT_TEMPR67[38] , \B_DOUT_TEMPR68[38] , 
        \B_DOUT_TEMPR69[38] , \B_DOUT_TEMPR70[38] , 
        \B_DOUT_TEMPR71[38] , \B_DOUT_TEMPR72[38] , 
        \B_DOUT_TEMPR73[38] , \B_DOUT_TEMPR74[38] , 
        \B_DOUT_TEMPR75[38] , \B_DOUT_TEMPR76[38] , 
        \B_DOUT_TEMPR77[38] , \B_DOUT_TEMPR78[38] , 
        \B_DOUT_TEMPR79[38] , \B_DOUT_TEMPR80[38] , 
        \B_DOUT_TEMPR81[38] , \B_DOUT_TEMPR82[38] , 
        \B_DOUT_TEMPR83[38] , \B_DOUT_TEMPR84[38] , 
        \B_DOUT_TEMPR85[38] , \B_DOUT_TEMPR86[38] , 
        \B_DOUT_TEMPR87[38] , \B_DOUT_TEMPR88[38] , 
        \B_DOUT_TEMPR89[38] , \B_DOUT_TEMPR90[38] , 
        \B_DOUT_TEMPR91[38] , \B_DOUT_TEMPR92[38] , 
        \B_DOUT_TEMPR93[38] , \B_DOUT_TEMPR94[38] , 
        \B_DOUT_TEMPR95[38] , \B_DOUT_TEMPR96[38] , 
        \B_DOUT_TEMPR97[38] , \B_DOUT_TEMPR98[38] , 
        \B_DOUT_TEMPR99[38] , \B_DOUT_TEMPR100[38] , 
        \B_DOUT_TEMPR101[38] , \B_DOUT_TEMPR102[38] , 
        \B_DOUT_TEMPR103[38] , \B_DOUT_TEMPR104[38] , 
        \B_DOUT_TEMPR105[38] , \B_DOUT_TEMPR106[38] , 
        \B_DOUT_TEMPR107[38] , \B_DOUT_TEMPR108[38] , 
        \B_DOUT_TEMPR109[38] , \B_DOUT_TEMPR110[38] , 
        \B_DOUT_TEMPR111[38] , \B_DOUT_TEMPR112[38] , 
        \B_DOUT_TEMPR113[38] , \B_DOUT_TEMPR114[38] , 
        \B_DOUT_TEMPR115[38] , \B_DOUT_TEMPR116[38] , 
        \B_DOUT_TEMPR117[38] , \B_DOUT_TEMPR118[38] , 
        \B_DOUT_TEMPR0[39] , \B_DOUT_TEMPR1[39] , \B_DOUT_TEMPR2[39] , 
        \B_DOUT_TEMPR3[39] , \B_DOUT_TEMPR4[39] , \B_DOUT_TEMPR5[39] , 
        \B_DOUT_TEMPR6[39] , \B_DOUT_TEMPR7[39] , \B_DOUT_TEMPR8[39] , 
        \B_DOUT_TEMPR9[39] , \B_DOUT_TEMPR10[39] , 
        \B_DOUT_TEMPR11[39] , \B_DOUT_TEMPR12[39] , 
        \B_DOUT_TEMPR13[39] , \B_DOUT_TEMPR14[39] , 
        \B_DOUT_TEMPR15[39] , \B_DOUT_TEMPR16[39] , 
        \B_DOUT_TEMPR17[39] , \B_DOUT_TEMPR18[39] , 
        \B_DOUT_TEMPR19[39] , \B_DOUT_TEMPR20[39] , 
        \B_DOUT_TEMPR21[39] , \B_DOUT_TEMPR22[39] , 
        \B_DOUT_TEMPR23[39] , \B_DOUT_TEMPR24[39] , 
        \B_DOUT_TEMPR25[39] , \B_DOUT_TEMPR26[39] , 
        \B_DOUT_TEMPR27[39] , \B_DOUT_TEMPR28[39] , 
        \B_DOUT_TEMPR29[39] , \B_DOUT_TEMPR30[39] , 
        \B_DOUT_TEMPR31[39] , \B_DOUT_TEMPR32[39] , 
        \B_DOUT_TEMPR33[39] , \B_DOUT_TEMPR34[39] , 
        \B_DOUT_TEMPR35[39] , \B_DOUT_TEMPR36[39] , 
        \B_DOUT_TEMPR37[39] , \B_DOUT_TEMPR38[39] , 
        \B_DOUT_TEMPR39[39] , \B_DOUT_TEMPR40[39] , 
        \B_DOUT_TEMPR41[39] , \B_DOUT_TEMPR42[39] , 
        \B_DOUT_TEMPR43[39] , \B_DOUT_TEMPR44[39] , 
        \B_DOUT_TEMPR45[39] , \B_DOUT_TEMPR46[39] , 
        \B_DOUT_TEMPR47[39] , \B_DOUT_TEMPR48[39] , 
        \B_DOUT_TEMPR49[39] , \B_DOUT_TEMPR50[39] , 
        \B_DOUT_TEMPR51[39] , \B_DOUT_TEMPR52[39] , 
        \B_DOUT_TEMPR53[39] , \B_DOUT_TEMPR54[39] , 
        \B_DOUT_TEMPR55[39] , \B_DOUT_TEMPR56[39] , 
        \B_DOUT_TEMPR57[39] , \B_DOUT_TEMPR58[39] , 
        \B_DOUT_TEMPR59[39] , \B_DOUT_TEMPR60[39] , 
        \B_DOUT_TEMPR61[39] , \B_DOUT_TEMPR62[39] , 
        \B_DOUT_TEMPR63[39] , \B_DOUT_TEMPR64[39] , 
        \B_DOUT_TEMPR65[39] , \B_DOUT_TEMPR66[39] , 
        \B_DOUT_TEMPR67[39] , \B_DOUT_TEMPR68[39] , 
        \B_DOUT_TEMPR69[39] , \B_DOUT_TEMPR70[39] , 
        \B_DOUT_TEMPR71[39] , \B_DOUT_TEMPR72[39] , 
        \B_DOUT_TEMPR73[39] , \B_DOUT_TEMPR74[39] , 
        \B_DOUT_TEMPR75[39] , \B_DOUT_TEMPR76[39] , 
        \B_DOUT_TEMPR77[39] , \B_DOUT_TEMPR78[39] , 
        \B_DOUT_TEMPR79[39] , \B_DOUT_TEMPR80[39] , 
        \B_DOUT_TEMPR81[39] , \B_DOUT_TEMPR82[39] , 
        \B_DOUT_TEMPR83[39] , \B_DOUT_TEMPR84[39] , 
        \B_DOUT_TEMPR85[39] , \B_DOUT_TEMPR86[39] , 
        \B_DOUT_TEMPR87[39] , \B_DOUT_TEMPR88[39] , 
        \B_DOUT_TEMPR89[39] , \B_DOUT_TEMPR90[39] , 
        \B_DOUT_TEMPR91[39] , \B_DOUT_TEMPR92[39] , 
        \B_DOUT_TEMPR93[39] , \B_DOUT_TEMPR94[39] , 
        \B_DOUT_TEMPR95[39] , \B_DOUT_TEMPR96[39] , 
        \B_DOUT_TEMPR97[39] , \B_DOUT_TEMPR98[39] , 
        \B_DOUT_TEMPR99[39] , \B_DOUT_TEMPR100[39] , 
        \B_DOUT_TEMPR101[39] , \B_DOUT_TEMPR102[39] , 
        \B_DOUT_TEMPR103[39] , \B_DOUT_TEMPR104[39] , 
        \B_DOUT_TEMPR105[39] , \B_DOUT_TEMPR106[39] , 
        \B_DOUT_TEMPR107[39] , \B_DOUT_TEMPR108[39] , 
        \B_DOUT_TEMPR109[39] , \B_DOUT_TEMPR110[39] , 
        \B_DOUT_TEMPR111[39] , \B_DOUT_TEMPR112[39] , 
        \B_DOUT_TEMPR113[39] , \B_DOUT_TEMPR114[39] , 
        \B_DOUT_TEMPR115[39] , \B_DOUT_TEMPR116[39] , 
        \B_DOUT_TEMPR117[39] , \B_DOUT_TEMPR118[39] , 
        \A_DOUT_TEMPR0[0] , \A_DOUT_TEMPR1[0] , \A_DOUT_TEMPR2[0] , 
        \A_DOUT_TEMPR3[0] , \A_DOUT_TEMPR4[0] , \A_DOUT_TEMPR5[0] , 
        \A_DOUT_TEMPR6[0] , \A_DOUT_TEMPR7[0] , \A_DOUT_TEMPR8[0] , 
        \A_DOUT_TEMPR9[0] , \A_DOUT_TEMPR10[0] , \A_DOUT_TEMPR11[0] , 
        \A_DOUT_TEMPR12[0] , \A_DOUT_TEMPR13[0] , \A_DOUT_TEMPR14[0] , 
        \A_DOUT_TEMPR15[0] , \A_DOUT_TEMPR16[0] , \A_DOUT_TEMPR17[0] , 
        \A_DOUT_TEMPR18[0] , \A_DOUT_TEMPR19[0] , \A_DOUT_TEMPR20[0] , 
        \A_DOUT_TEMPR21[0] , \A_DOUT_TEMPR22[0] , \A_DOUT_TEMPR23[0] , 
        \A_DOUT_TEMPR24[0] , \A_DOUT_TEMPR25[0] , \A_DOUT_TEMPR26[0] , 
        \A_DOUT_TEMPR27[0] , \A_DOUT_TEMPR28[0] , \A_DOUT_TEMPR29[0] , 
        \A_DOUT_TEMPR30[0] , \A_DOUT_TEMPR31[0] , \A_DOUT_TEMPR32[0] , 
        \A_DOUT_TEMPR33[0] , \A_DOUT_TEMPR34[0] , \A_DOUT_TEMPR35[0] , 
        \A_DOUT_TEMPR36[0] , \A_DOUT_TEMPR37[0] , \A_DOUT_TEMPR38[0] , 
        \A_DOUT_TEMPR39[0] , \A_DOUT_TEMPR40[0] , \A_DOUT_TEMPR41[0] , 
        \A_DOUT_TEMPR42[0] , \A_DOUT_TEMPR43[0] , \A_DOUT_TEMPR44[0] , 
        \A_DOUT_TEMPR45[0] , \A_DOUT_TEMPR46[0] , \A_DOUT_TEMPR47[0] , 
        \A_DOUT_TEMPR48[0] , \A_DOUT_TEMPR49[0] , \A_DOUT_TEMPR50[0] , 
        \A_DOUT_TEMPR51[0] , \A_DOUT_TEMPR52[0] , \A_DOUT_TEMPR53[0] , 
        \A_DOUT_TEMPR54[0] , \A_DOUT_TEMPR55[0] , \A_DOUT_TEMPR56[0] , 
        \A_DOUT_TEMPR57[0] , \A_DOUT_TEMPR58[0] , \A_DOUT_TEMPR59[0] , 
        \A_DOUT_TEMPR60[0] , \A_DOUT_TEMPR61[0] , \A_DOUT_TEMPR62[0] , 
        \A_DOUT_TEMPR63[0] , \A_DOUT_TEMPR64[0] , \A_DOUT_TEMPR65[0] , 
        \A_DOUT_TEMPR66[0] , \A_DOUT_TEMPR67[0] , \A_DOUT_TEMPR68[0] , 
        \A_DOUT_TEMPR69[0] , \A_DOUT_TEMPR70[0] , \A_DOUT_TEMPR71[0] , 
        \A_DOUT_TEMPR72[0] , \A_DOUT_TEMPR73[0] , \A_DOUT_TEMPR74[0] , 
        \A_DOUT_TEMPR75[0] , \A_DOUT_TEMPR76[0] , \A_DOUT_TEMPR77[0] , 
        \A_DOUT_TEMPR78[0] , \A_DOUT_TEMPR79[0] , \A_DOUT_TEMPR80[0] , 
        \A_DOUT_TEMPR81[0] , \A_DOUT_TEMPR82[0] , \A_DOUT_TEMPR83[0] , 
        \A_DOUT_TEMPR84[0] , \A_DOUT_TEMPR85[0] , \A_DOUT_TEMPR86[0] , 
        \A_DOUT_TEMPR87[0] , \A_DOUT_TEMPR88[0] , \A_DOUT_TEMPR89[0] , 
        \A_DOUT_TEMPR90[0] , \A_DOUT_TEMPR91[0] , \A_DOUT_TEMPR92[0] , 
        \A_DOUT_TEMPR93[0] , \A_DOUT_TEMPR94[0] , \A_DOUT_TEMPR95[0] , 
        \A_DOUT_TEMPR96[0] , \A_DOUT_TEMPR97[0] , \A_DOUT_TEMPR98[0] , 
        \A_DOUT_TEMPR99[0] , \A_DOUT_TEMPR100[0] , 
        \A_DOUT_TEMPR101[0] , \A_DOUT_TEMPR102[0] , 
        \A_DOUT_TEMPR103[0] , \A_DOUT_TEMPR104[0] , 
        \A_DOUT_TEMPR105[0] , \A_DOUT_TEMPR106[0] , 
        \A_DOUT_TEMPR107[0] , \A_DOUT_TEMPR108[0] , 
        \A_DOUT_TEMPR109[0] , \A_DOUT_TEMPR110[0] , 
        \A_DOUT_TEMPR111[0] , \A_DOUT_TEMPR112[0] , 
        \A_DOUT_TEMPR113[0] , \A_DOUT_TEMPR114[0] , 
        \A_DOUT_TEMPR115[0] , \A_DOUT_TEMPR116[0] , 
        \A_DOUT_TEMPR117[0] , \A_DOUT_TEMPR118[0] , \A_DOUT_TEMPR0[1] , 
        \A_DOUT_TEMPR1[1] , \A_DOUT_TEMPR2[1] , \A_DOUT_TEMPR3[1] , 
        \A_DOUT_TEMPR4[1] , \A_DOUT_TEMPR5[1] , \A_DOUT_TEMPR6[1] , 
        \A_DOUT_TEMPR7[1] , \A_DOUT_TEMPR8[1] , \A_DOUT_TEMPR9[1] , 
        \A_DOUT_TEMPR10[1] , \A_DOUT_TEMPR11[1] , \A_DOUT_TEMPR12[1] , 
        \A_DOUT_TEMPR13[1] , \A_DOUT_TEMPR14[1] , \A_DOUT_TEMPR15[1] , 
        \A_DOUT_TEMPR16[1] , \A_DOUT_TEMPR17[1] , \A_DOUT_TEMPR18[1] , 
        \A_DOUT_TEMPR19[1] , \A_DOUT_TEMPR20[1] , \A_DOUT_TEMPR21[1] , 
        \A_DOUT_TEMPR22[1] , \A_DOUT_TEMPR23[1] , \A_DOUT_TEMPR24[1] , 
        \A_DOUT_TEMPR25[1] , \A_DOUT_TEMPR26[1] , \A_DOUT_TEMPR27[1] , 
        \A_DOUT_TEMPR28[1] , \A_DOUT_TEMPR29[1] , \A_DOUT_TEMPR30[1] , 
        \A_DOUT_TEMPR31[1] , \A_DOUT_TEMPR32[1] , \A_DOUT_TEMPR33[1] , 
        \A_DOUT_TEMPR34[1] , \A_DOUT_TEMPR35[1] , \A_DOUT_TEMPR36[1] , 
        \A_DOUT_TEMPR37[1] , \A_DOUT_TEMPR38[1] , \A_DOUT_TEMPR39[1] , 
        \A_DOUT_TEMPR40[1] , \A_DOUT_TEMPR41[1] , \A_DOUT_TEMPR42[1] , 
        \A_DOUT_TEMPR43[1] , \A_DOUT_TEMPR44[1] , \A_DOUT_TEMPR45[1] , 
        \A_DOUT_TEMPR46[1] , \A_DOUT_TEMPR47[1] , \A_DOUT_TEMPR48[1] , 
        \A_DOUT_TEMPR49[1] , \A_DOUT_TEMPR50[1] , \A_DOUT_TEMPR51[1] , 
        \A_DOUT_TEMPR52[1] , \A_DOUT_TEMPR53[1] , \A_DOUT_TEMPR54[1] , 
        \A_DOUT_TEMPR55[1] , \A_DOUT_TEMPR56[1] , \A_DOUT_TEMPR57[1] , 
        \A_DOUT_TEMPR58[1] , \A_DOUT_TEMPR59[1] , \A_DOUT_TEMPR60[1] , 
        \A_DOUT_TEMPR61[1] , \A_DOUT_TEMPR62[1] , \A_DOUT_TEMPR63[1] , 
        \A_DOUT_TEMPR64[1] , \A_DOUT_TEMPR65[1] , \A_DOUT_TEMPR66[1] , 
        \A_DOUT_TEMPR67[1] , \A_DOUT_TEMPR68[1] , \A_DOUT_TEMPR69[1] , 
        \A_DOUT_TEMPR70[1] , \A_DOUT_TEMPR71[1] , \A_DOUT_TEMPR72[1] , 
        \A_DOUT_TEMPR73[1] , \A_DOUT_TEMPR74[1] , \A_DOUT_TEMPR75[1] , 
        \A_DOUT_TEMPR76[1] , \A_DOUT_TEMPR77[1] , \A_DOUT_TEMPR78[1] , 
        \A_DOUT_TEMPR79[1] , \A_DOUT_TEMPR80[1] , \A_DOUT_TEMPR81[1] , 
        \A_DOUT_TEMPR82[1] , \A_DOUT_TEMPR83[1] , \A_DOUT_TEMPR84[1] , 
        \A_DOUT_TEMPR85[1] , \A_DOUT_TEMPR86[1] , \A_DOUT_TEMPR87[1] , 
        \A_DOUT_TEMPR88[1] , \A_DOUT_TEMPR89[1] , \A_DOUT_TEMPR90[1] , 
        \A_DOUT_TEMPR91[1] , \A_DOUT_TEMPR92[1] , \A_DOUT_TEMPR93[1] , 
        \A_DOUT_TEMPR94[1] , \A_DOUT_TEMPR95[1] , \A_DOUT_TEMPR96[1] , 
        \A_DOUT_TEMPR97[1] , \A_DOUT_TEMPR98[1] , \A_DOUT_TEMPR99[1] , 
        \A_DOUT_TEMPR100[1] , \A_DOUT_TEMPR101[1] , 
        \A_DOUT_TEMPR102[1] , \A_DOUT_TEMPR103[1] , 
        \A_DOUT_TEMPR104[1] , \A_DOUT_TEMPR105[1] , 
        \A_DOUT_TEMPR106[1] , \A_DOUT_TEMPR107[1] , 
        \A_DOUT_TEMPR108[1] , \A_DOUT_TEMPR109[1] , 
        \A_DOUT_TEMPR110[1] , \A_DOUT_TEMPR111[1] , 
        \A_DOUT_TEMPR112[1] , \A_DOUT_TEMPR113[1] , 
        \A_DOUT_TEMPR114[1] , \A_DOUT_TEMPR115[1] , 
        \A_DOUT_TEMPR116[1] , \A_DOUT_TEMPR117[1] , 
        \A_DOUT_TEMPR118[1] , \A_DOUT_TEMPR0[2] , \A_DOUT_TEMPR1[2] , 
        \A_DOUT_TEMPR2[2] , \A_DOUT_TEMPR3[2] , \A_DOUT_TEMPR4[2] , 
        \A_DOUT_TEMPR5[2] , \A_DOUT_TEMPR6[2] , \A_DOUT_TEMPR7[2] , 
        \A_DOUT_TEMPR8[2] , \A_DOUT_TEMPR9[2] , \A_DOUT_TEMPR10[2] , 
        \A_DOUT_TEMPR11[2] , \A_DOUT_TEMPR12[2] , \A_DOUT_TEMPR13[2] , 
        \A_DOUT_TEMPR14[2] , \A_DOUT_TEMPR15[2] , \A_DOUT_TEMPR16[2] , 
        \A_DOUT_TEMPR17[2] , \A_DOUT_TEMPR18[2] , \A_DOUT_TEMPR19[2] , 
        \A_DOUT_TEMPR20[2] , \A_DOUT_TEMPR21[2] , \A_DOUT_TEMPR22[2] , 
        \A_DOUT_TEMPR23[2] , \A_DOUT_TEMPR24[2] , \A_DOUT_TEMPR25[2] , 
        \A_DOUT_TEMPR26[2] , \A_DOUT_TEMPR27[2] , \A_DOUT_TEMPR28[2] , 
        \A_DOUT_TEMPR29[2] , \A_DOUT_TEMPR30[2] , \A_DOUT_TEMPR31[2] , 
        \A_DOUT_TEMPR32[2] , \A_DOUT_TEMPR33[2] , \A_DOUT_TEMPR34[2] , 
        \A_DOUT_TEMPR35[2] , \A_DOUT_TEMPR36[2] , \A_DOUT_TEMPR37[2] , 
        \A_DOUT_TEMPR38[2] , \A_DOUT_TEMPR39[2] , \A_DOUT_TEMPR40[2] , 
        \A_DOUT_TEMPR41[2] , \A_DOUT_TEMPR42[2] , \A_DOUT_TEMPR43[2] , 
        \A_DOUT_TEMPR44[2] , \A_DOUT_TEMPR45[2] , \A_DOUT_TEMPR46[2] , 
        \A_DOUT_TEMPR47[2] , \A_DOUT_TEMPR48[2] , \A_DOUT_TEMPR49[2] , 
        \A_DOUT_TEMPR50[2] , \A_DOUT_TEMPR51[2] , \A_DOUT_TEMPR52[2] , 
        \A_DOUT_TEMPR53[2] , \A_DOUT_TEMPR54[2] , \A_DOUT_TEMPR55[2] , 
        \A_DOUT_TEMPR56[2] , \A_DOUT_TEMPR57[2] , \A_DOUT_TEMPR58[2] , 
        \A_DOUT_TEMPR59[2] , \A_DOUT_TEMPR60[2] , \A_DOUT_TEMPR61[2] , 
        \A_DOUT_TEMPR62[2] , \A_DOUT_TEMPR63[2] , \A_DOUT_TEMPR64[2] , 
        \A_DOUT_TEMPR65[2] , \A_DOUT_TEMPR66[2] , \A_DOUT_TEMPR67[2] , 
        \A_DOUT_TEMPR68[2] , \A_DOUT_TEMPR69[2] , \A_DOUT_TEMPR70[2] , 
        \A_DOUT_TEMPR71[2] , \A_DOUT_TEMPR72[2] , \A_DOUT_TEMPR73[2] , 
        \A_DOUT_TEMPR74[2] , \A_DOUT_TEMPR75[2] , \A_DOUT_TEMPR76[2] , 
        \A_DOUT_TEMPR77[2] , \A_DOUT_TEMPR78[2] , \A_DOUT_TEMPR79[2] , 
        \A_DOUT_TEMPR80[2] , \A_DOUT_TEMPR81[2] , \A_DOUT_TEMPR82[2] , 
        \A_DOUT_TEMPR83[2] , \A_DOUT_TEMPR84[2] , \A_DOUT_TEMPR85[2] , 
        \A_DOUT_TEMPR86[2] , \A_DOUT_TEMPR87[2] , \A_DOUT_TEMPR88[2] , 
        \A_DOUT_TEMPR89[2] , \A_DOUT_TEMPR90[2] , \A_DOUT_TEMPR91[2] , 
        \A_DOUT_TEMPR92[2] , \A_DOUT_TEMPR93[2] , \A_DOUT_TEMPR94[2] , 
        \A_DOUT_TEMPR95[2] , \A_DOUT_TEMPR96[2] , \A_DOUT_TEMPR97[2] , 
        \A_DOUT_TEMPR98[2] , \A_DOUT_TEMPR99[2] , \A_DOUT_TEMPR100[2] , 
        \A_DOUT_TEMPR101[2] , \A_DOUT_TEMPR102[2] , 
        \A_DOUT_TEMPR103[2] , \A_DOUT_TEMPR104[2] , 
        \A_DOUT_TEMPR105[2] , \A_DOUT_TEMPR106[2] , 
        \A_DOUT_TEMPR107[2] , \A_DOUT_TEMPR108[2] , 
        \A_DOUT_TEMPR109[2] , \A_DOUT_TEMPR110[2] , 
        \A_DOUT_TEMPR111[2] , \A_DOUT_TEMPR112[2] , 
        \A_DOUT_TEMPR113[2] , \A_DOUT_TEMPR114[2] , 
        \A_DOUT_TEMPR115[2] , \A_DOUT_TEMPR116[2] , 
        \A_DOUT_TEMPR117[2] , \A_DOUT_TEMPR118[2] , \A_DOUT_TEMPR0[3] , 
        \A_DOUT_TEMPR1[3] , \A_DOUT_TEMPR2[3] , \A_DOUT_TEMPR3[3] , 
        \A_DOUT_TEMPR4[3] , \A_DOUT_TEMPR5[3] , \A_DOUT_TEMPR6[3] , 
        \A_DOUT_TEMPR7[3] , \A_DOUT_TEMPR8[3] , \A_DOUT_TEMPR9[3] , 
        \A_DOUT_TEMPR10[3] , \A_DOUT_TEMPR11[3] , \A_DOUT_TEMPR12[3] , 
        \A_DOUT_TEMPR13[3] , \A_DOUT_TEMPR14[3] , \A_DOUT_TEMPR15[3] , 
        \A_DOUT_TEMPR16[3] , \A_DOUT_TEMPR17[3] , \A_DOUT_TEMPR18[3] , 
        \A_DOUT_TEMPR19[3] , \A_DOUT_TEMPR20[3] , \A_DOUT_TEMPR21[3] , 
        \A_DOUT_TEMPR22[3] , \A_DOUT_TEMPR23[3] , \A_DOUT_TEMPR24[3] , 
        \A_DOUT_TEMPR25[3] , \A_DOUT_TEMPR26[3] , \A_DOUT_TEMPR27[3] , 
        \A_DOUT_TEMPR28[3] , \A_DOUT_TEMPR29[3] , \A_DOUT_TEMPR30[3] , 
        \A_DOUT_TEMPR31[3] , \A_DOUT_TEMPR32[3] , \A_DOUT_TEMPR33[3] , 
        \A_DOUT_TEMPR34[3] , \A_DOUT_TEMPR35[3] , \A_DOUT_TEMPR36[3] , 
        \A_DOUT_TEMPR37[3] , \A_DOUT_TEMPR38[3] , \A_DOUT_TEMPR39[3] , 
        \A_DOUT_TEMPR40[3] , \A_DOUT_TEMPR41[3] , \A_DOUT_TEMPR42[3] , 
        \A_DOUT_TEMPR43[3] , \A_DOUT_TEMPR44[3] , \A_DOUT_TEMPR45[3] , 
        \A_DOUT_TEMPR46[3] , \A_DOUT_TEMPR47[3] , \A_DOUT_TEMPR48[3] , 
        \A_DOUT_TEMPR49[3] , \A_DOUT_TEMPR50[3] , \A_DOUT_TEMPR51[3] , 
        \A_DOUT_TEMPR52[3] , \A_DOUT_TEMPR53[3] , \A_DOUT_TEMPR54[3] , 
        \A_DOUT_TEMPR55[3] , \A_DOUT_TEMPR56[3] , \A_DOUT_TEMPR57[3] , 
        \A_DOUT_TEMPR58[3] , \A_DOUT_TEMPR59[3] , \A_DOUT_TEMPR60[3] , 
        \A_DOUT_TEMPR61[3] , \A_DOUT_TEMPR62[3] , \A_DOUT_TEMPR63[3] , 
        \A_DOUT_TEMPR64[3] , \A_DOUT_TEMPR65[3] , \A_DOUT_TEMPR66[3] , 
        \A_DOUT_TEMPR67[3] , \A_DOUT_TEMPR68[3] , \A_DOUT_TEMPR69[3] , 
        \A_DOUT_TEMPR70[3] , \A_DOUT_TEMPR71[3] , \A_DOUT_TEMPR72[3] , 
        \A_DOUT_TEMPR73[3] , \A_DOUT_TEMPR74[3] , \A_DOUT_TEMPR75[3] , 
        \A_DOUT_TEMPR76[3] , \A_DOUT_TEMPR77[3] , \A_DOUT_TEMPR78[3] , 
        \A_DOUT_TEMPR79[3] , \A_DOUT_TEMPR80[3] , \A_DOUT_TEMPR81[3] , 
        \A_DOUT_TEMPR82[3] , \A_DOUT_TEMPR83[3] , \A_DOUT_TEMPR84[3] , 
        \A_DOUT_TEMPR85[3] , \A_DOUT_TEMPR86[3] , \A_DOUT_TEMPR87[3] , 
        \A_DOUT_TEMPR88[3] , \A_DOUT_TEMPR89[3] , \A_DOUT_TEMPR90[3] , 
        \A_DOUT_TEMPR91[3] , \A_DOUT_TEMPR92[3] , \A_DOUT_TEMPR93[3] , 
        \A_DOUT_TEMPR94[3] , \A_DOUT_TEMPR95[3] , \A_DOUT_TEMPR96[3] , 
        \A_DOUT_TEMPR97[3] , \A_DOUT_TEMPR98[3] , \A_DOUT_TEMPR99[3] , 
        \A_DOUT_TEMPR100[3] , \A_DOUT_TEMPR101[3] , 
        \A_DOUT_TEMPR102[3] , \A_DOUT_TEMPR103[3] , 
        \A_DOUT_TEMPR104[3] , \A_DOUT_TEMPR105[3] , 
        \A_DOUT_TEMPR106[3] , \A_DOUT_TEMPR107[3] , 
        \A_DOUT_TEMPR108[3] , \A_DOUT_TEMPR109[3] , 
        \A_DOUT_TEMPR110[3] , \A_DOUT_TEMPR111[3] , 
        \A_DOUT_TEMPR112[3] , \A_DOUT_TEMPR113[3] , 
        \A_DOUT_TEMPR114[3] , \A_DOUT_TEMPR115[3] , 
        \A_DOUT_TEMPR116[3] , \A_DOUT_TEMPR117[3] , 
        \A_DOUT_TEMPR118[3] , \A_DOUT_TEMPR0[4] , \A_DOUT_TEMPR1[4] , 
        \A_DOUT_TEMPR2[4] , \A_DOUT_TEMPR3[4] , \A_DOUT_TEMPR4[4] , 
        \A_DOUT_TEMPR5[4] , \A_DOUT_TEMPR6[4] , \A_DOUT_TEMPR7[4] , 
        \A_DOUT_TEMPR8[4] , \A_DOUT_TEMPR9[4] , \A_DOUT_TEMPR10[4] , 
        \A_DOUT_TEMPR11[4] , \A_DOUT_TEMPR12[4] , \A_DOUT_TEMPR13[4] , 
        \A_DOUT_TEMPR14[4] , \A_DOUT_TEMPR15[4] , \A_DOUT_TEMPR16[4] , 
        \A_DOUT_TEMPR17[4] , \A_DOUT_TEMPR18[4] , \A_DOUT_TEMPR19[4] , 
        \A_DOUT_TEMPR20[4] , \A_DOUT_TEMPR21[4] , \A_DOUT_TEMPR22[4] , 
        \A_DOUT_TEMPR23[4] , \A_DOUT_TEMPR24[4] , \A_DOUT_TEMPR25[4] , 
        \A_DOUT_TEMPR26[4] , \A_DOUT_TEMPR27[4] , \A_DOUT_TEMPR28[4] , 
        \A_DOUT_TEMPR29[4] , \A_DOUT_TEMPR30[4] , \A_DOUT_TEMPR31[4] , 
        \A_DOUT_TEMPR32[4] , \A_DOUT_TEMPR33[4] , \A_DOUT_TEMPR34[4] , 
        \A_DOUT_TEMPR35[4] , \A_DOUT_TEMPR36[4] , \A_DOUT_TEMPR37[4] , 
        \A_DOUT_TEMPR38[4] , \A_DOUT_TEMPR39[4] , \A_DOUT_TEMPR40[4] , 
        \A_DOUT_TEMPR41[4] , \A_DOUT_TEMPR42[4] , \A_DOUT_TEMPR43[4] , 
        \A_DOUT_TEMPR44[4] , \A_DOUT_TEMPR45[4] , \A_DOUT_TEMPR46[4] , 
        \A_DOUT_TEMPR47[4] , \A_DOUT_TEMPR48[4] , \A_DOUT_TEMPR49[4] , 
        \A_DOUT_TEMPR50[4] , \A_DOUT_TEMPR51[4] , \A_DOUT_TEMPR52[4] , 
        \A_DOUT_TEMPR53[4] , \A_DOUT_TEMPR54[4] , \A_DOUT_TEMPR55[4] , 
        \A_DOUT_TEMPR56[4] , \A_DOUT_TEMPR57[4] , \A_DOUT_TEMPR58[4] , 
        \A_DOUT_TEMPR59[4] , \A_DOUT_TEMPR60[4] , \A_DOUT_TEMPR61[4] , 
        \A_DOUT_TEMPR62[4] , \A_DOUT_TEMPR63[4] , \A_DOUT_TEMPR64[4] , 
        \A_DOUT_TEMPR65[4] , \A_DOUT_TEMPR66[4] , \A_DOUT_TEMPR67[4] , 
        \A_DOUT_TEMPR68[4] , \A_DOUT_TEMPR69[4] , \A_DOUT_TEMPR70[4] , 
        \A_DOUT_TEMPR71[4] , \A_DOUT_TEMPR72[4] , \A_DOUT_TEMPR73[4] , 
        \A_DOUT_TEMPR74[4] , \A_DOUT_TEMPR75[4] , \A_DOUT_TEMPR76[4] , 
        \A_DOUT_TEMPR77[4] , \A_DOUT_TEMPR78[4] , \A_DOUT_TEMPR79[4] , 
        \A_DOUT_TEMPR80[4] , \A_DOUT_TEMPR81[4] , \A_DOUT_TEMPR82[4] , 
        \A_DOUT_TEMPR83[4] , \A_DOUT_TEMPR84[4] , \A_DOUT_TEMPR85[4] , 
        \A_DOUT_TEMPR86[4] , \A_DOUT_TEMPR87[4] , \A_DOUT_TEMPR88[4] , 
        \A_DOUT_TEMPR89[4] , \A_DOUT_TEMPR90[4] , \A_DOUT_TEMPR91[4] , 
        \A_DOUT_TEMPR92[4] , \A_DOUT_TEMPR93[4] , \A_DOUT_TEMPR94[4] , 
        \A_DOUT_TEMPR95[4] , \A_DOUT_TEMPR96[4] , \A_DOUT_TEMPR97[4] , 
        \A_DOUT_TEMPR98[4] , \A_DOUT_TEMPR99[4] , \A_DOUT_TEMPR100[4] , 
        \A_DOUT_TEMPR101[4] , \A_DOUT_TEMPR102[4] , 
        \A_DOUT_TEMPR103[4] , \A_DOUT_TEMPR104[4] , 
        \A_DOUT_TEMPR105[4] , \A_DOUT_TEMPR106[4] , 
        \A_DOUT_TEMPR107[4] , \A_DOUT_TEMPR108[4] , 
        \A_DOUT_TEMPR109[4] , \A_DOUT_TEMPR110[4] , 
        \A_DOUT_TEMPR111[4] , \A_DOUT_TEMPR112[4] , 
        \A_DOUT_TEMPR113[4] , \A_DOUT_TEMPR114[4] , 
        \A_DOUT_TEMPR115[4] , \A_DOUT_TEMPR116[4] , 
        \A_DOUT_TEMPR117[4] , \A_DOUT_TEMPR118[4] , \A_DOUT_TEMPR0[5] , 
        \A_DOUT_TEMPR1[5] , \A_DOUT_TEMPR2[5] , \A_DOUT_TEMPR3[5] , 
        \A_DOUT_TEMPR4[5] , \A_DOUT_TEMPR5[5] , \A_DOUT_TEMPR6[5] , 
        \A_DOUT_TEMPR7[5] , \A_DOUT_TEMPR8[5] , \A_DOUT_TEMPR9[5] , 
        \A_DOUT_TEMPR10[5] , \A_DOUT_TEMPR11[5] , \A_DOUT_TEMPR12[5] , 
        \A_DOUT_TEMPR13[5] , \A_DOUT_TEMPR14[5] , \A_DOUT_TEMPR15[5] , 
        \A_DOUT_TEMPR16[5] , \A_DOUT_TEMPR17[5] , \A_DOUT_TEMPR18[5] , 
        \A_DOUT_TEMPR19[5] , \A_DOUT_TEMPR20[5] , \A_DOUT_TEMPR21[5] , 
        \A_DOUT_TEMPR22[5] , \A_DOUT_TEMPR23[5] , \A_DOUT_TEMPR24[5] , 
        \A_DOUT_TEMPR25[5] , \A_DOUT_TEMPR26[5] , \A_DOUT_TEMPR27[5] , 
        \A_DOUT_TEMPR28[5] , \A_DOUT_TEMPR29[5] , \A_DOUT_TEMPR30[5] , 
        \A_DOUT_TEMPR31[5] , \A_DOUT_TEMPR32[5] , \A_DOUT_TEMPR33[5] , 
        \A_DOUT_TEMPR34[5] , \A_DOUT_TEMPR35[5] , \A_DOUT_TEMPR36[5] , 
        \A_DOUT_TEMPR37[5] , \A_DOUT_TEMPR38[5] , \A_DOUT_TEMPR39[5] , 
        \A_DOUT_TEMPR40[5] , \A_DOUT_TEMPR41[5] , \A_DOUT_TEMPR42[5] , 
        \A_DOUT_TEMPR43[5] , \A_DOUT_TEMPR44[5] , \A_DOUT_TEMPR45[5] , 
        \A_DOUT_TEMPR46[5] , \A_DOUT_TEMPR47[5] , \A_DOUT_TEMPR48[5] , 
        \A_DOUT_TEMPR49[5] , \A_DOUT_TEMPR50[5] , \A_DOUT_TEMPR51[5] , 
        \A_DOUT_TEMPR52[5] , \A_DOUT_TEMPR53[5] , \A_DOUT_TEMPR54[5] , 
        \A_DOUT_TEMPR55[5] , \A_DOUT_TEMPR56[5] , \A_DOUT_TEMPR57[5] , 
        \A_DOUT_TEMPR58[5] , \A_DOUT_TEMPR59[5] , \A_DOUT_TEMPR60[5] , 
        \A_DOUT_TEMPR61[5] , \A_DOUT_TEMPR62[5] , \A_DOUT_TEMPR63[5] , 
        \A_DOUT_TEMPR64[5] , \A_DOUT_TEMPR65[5] , \A_DOUT_TEMPR66[5] , 
        \A_DOUT_TEMPR67[5] , \A_DOUT_TEMPR68[5] , \A_DOUT_TEMPR69[5] , 
        \A_DOUT_TEMPR70[5] , \A_DOUT_TEMPR71[5] , \A_DOUT_TEMPR72[5] , 
        \A_DOUT_TEMPR73[5] , \A_DOUT_TEMPR74[5] , \A_DOUT_TEMPR75[5] , 
        \A_DOUT_TEMPR76[5] , \A_DOUT_TEMPR77[5] , \A_DOUT_TEMPR78[5] , 
        \A_DOUT_TEMPR79[5] , \A_DOUT_TEMPR80[5] , \A_DOUT_TEMPR81[5] , 
        \A_DOUT_TEMPR82[5] , \A_DOUT_TEMPR83[5] , \A_DOUT_TEMPR84[5] , 
        \A_DOUT_TEMPR85[5] , \A_DOUT_TEMPR86[5] , \A_DOUT_TEMPR87[5] , 
        \A_DOUT_TEMPR88[5] , \A_DOUT_TEMPR89[5] , \A_DOUT_TEMPR90[5] , 
        \A_DOUT_TEMPR91[5] , \A_DOUT_TEMPR92[5] , \A_DOUT_TEMPR93[5] , 
        \A_DOUT_TEMPR94[5] , \A_DOUT_TEMPR95[5] , \A_DOUT_TEMPR96[5] , 
        \A_DOUT_TEMPR97[5] , \A_DOUT_TEMPR98[5] , \A_DOUT_TEMPR99[5] , 
        \A_DOUT_TEMPR100[5] , \A_DOUT_TEMPR101[5] , 
        \A_DOUT_TEMPR102[5] , \A_DOUT_TEMPR103[5] , 
        \A_DOUT_TEMPR104[5] , \A_DOUT_TEMPR105[5] , 
        \A_DOUT_TEMPR106[5] , \A_DOUT_TEMPR107[5] , 
        \A_DOUT_TEMPR108[5] , \A_DOUT_TEMPR109[5] , 
        \A_DOUT_TEMPR110[5] , \A_DOUT_TEMPR111[5] , 
        \A_DOUT_TEMPR112[5] , \A_DOUT_TEMPR113[5] , 
        \A_DOUT_TEMPR114[5] , \A_DOUT_TEMPR115[5] , 
        \A_DOUT_TEMPR116[5] , \A_DOUT_TEMPR117[5] , 
        \A_DOUT_TEMPR118[5] , \A_DOUT_TEMPR0[6] , \A_DOUT_TEMPR1[6] , 
        \A_DOUT_TEMPR2[6] , \A_DOUT_TEMPR3[6] , \A_DOUT_TEMPR4[6] , 
        \A_DOUT_TEMPR5[6] , \A_DOUT_TEMPR6[6] , \A_DOUT_TEMPR7[6] , 
        \A_DOUT_TEMPR8[6] , \A_DOUT_TEMPR9[6] , \A_DOUT_TEMPR10[6] , 
        \A_DOUT_TEMPR11[6] , \A_DOUT_TEMPR12[6] , \A_DOUT_TEMPR13[6] , 
        \A_DOUT_TEMPR14[6] , \A_DOUT_TEMPR15[6] , \A_DOUT_TEMPR16[6] , 
        \A_DOUT_TEMPR17[6] , \A_DOUT_TEMPR18[6] , \A_DOUT_TEMPR19[6] , 
        \A_DOUT_TEMPR20[6] , \A_DOUT_TEMPR21[6] , \A_DOUT_TEMPR22[6] , 
        \A_DOUT_TEMPR23[6] , \A_DOUT_TEMPR24[6] , \A_DOUT_TEMPR25[6] , 
        \A_DOUT_TEMPR26[6] , \A_DOUT_TEMPR27[6] , \A_DOUT_TEMPR28[6] , 
        \A_DOUT_TEMPR29[6] , \A_DOUT_TEMPR30[6] , \A_DOUT_TEMPR31[6] , 
        \A_DOUT_TEMPR32[6] , \A_DOUT_TEMPR33[6] , \A_DOUT_TEMPR34[6] , 
        \A_DOUT_TEMPR35[6] , \A_DOUT_TEMPR36[6] , \A_DOUT_TEMPR37[6] , 
        \A_DOUT_TEMPR38[6] , \A_DOUT_TEMPR39[6] , \A_DOUT_TEMPR40[6] , 
        \A_DOUT_TEMPR41[6] , \A_DOUT_TEMPR42[6] , \A_DOUT_TEMPR43[6] , 
        \A_DOUT_TEMPR44[6] , \A_DOUT_TEMPR45[6] , \A_DOUT_TEMPR46[6] , 
        \A_DOUT_TEMPR47[6] , \A_DOUT_TEMPR48[6] , \A_DOUT_TEMPR49[6] , 
        \A_DOUT_TEMPR50[6] , \A_DOUT_TEMPR51[6] , \A_DOUT_TEMPR52[6] , 
        \A_DOUT_TEMPR53[6] , \A_DOUT_TEMPR54[6] , \A_DOUT_TEMPR55[6] , 
        \A_DOUT_TEMPR56[6] , \A_DOUT_TEMPR57[6] , \A_DOUT_TEMPR58[6] , 
        \A_DOUT_TEMPR59[6] , \A_DOUT_TEMPR60[6] , \A_DOUT_TEMPR61[6] , 
        \A_DOUT_TEMPR62[6] , \A_DOUT_TEMPR63[6] , \A_DOUT_TEMPR64[6] , 
        \A_DOUT_TEMPR65[6] , \A_DOUT_TEMPR66[6] , \A_DOUT_TEMPR67[6] , 
        \A_DOUT_TEMPR68[6] , \A_DOUT_TEMPR69[6] , \A_DOUT_TEMPR70[6] , 
        \A_DOUT_TEMPR71[6] , \A_DOUT_TEMPR72[6] , \A_DOUT_TEMPR73[6] , 
        \A_DOUT_TEMPR74[6] , \A_DOUT_TEMPR75[6] , \A_DOUT_TEMPR76[6] , 
        \A_DOUT_TEMPR77[6] , \A_DOUT_TEMPR78[6] , \A_DOUT_TEMPR79[6] , 
        \A_DOUT_TEMPR80[6] , \A_DOUT_TEMPR81[6] , \A_DOUT_TEMPR82[6] , 
        \A_DOUT_TEMPR83[6] , \A_DOUT_TEMPR84[6] , \A_DOUT_TEMPR85[6] , 
        \A_DOUT_TEMPR86[6] , \A_DOUT_TEMPR87[6] , \A_DOUT_TEMPR88[6] , 
        \A_DOUT_TEMPR89[6] , \A_DOUT_TEMPR90[6] , \A_DOUT_TEMPR91[6] , 
        \A_DOUT_TEMPR92[6] , \A_DOUT_TEMPR93[6] , \A_DOUT_TEMPR94[6] , 
        \A_DOUT_TEMPR95[6] , \A_DOUT_TEMPR96[6] , \A_DOUT_TEMPR97[6] , 
        \A_DOUT_TEMPR98[6] , \A_DOUT_TEMPR99[6] , \A_DOUT_TEMPR100[6] , 
        \A_DOUT_TEMPR101[6] , \A_DOUT_TEMPR102[6] , 
        \A_DOUT_TEMPR103[6] , \A_DOUT_TEMPR104[6] , 
        \A_DOUT_TEMPR105[6] , \A_DOUT_TEMPR106[6] , 
        \A_DOUT_TEMPR107[6] , \A_DOUT_TEMPR108[6] , 
        \A_DOUT_TEMPR109[6] , \A_DOUT_TEMPR110[6] , 
        \A_DOUT_TEMPR111[6] , \A_DOUT_TEMPR112[6] , 
        \A_DOUT_TEMPR113[6] , \A_DOUT_TEMPR114[6] , 
        \A_DOUT_TEMPR115[6] , \A_DOUT_TEMPR116[6] , 
        \A_DOUT_TEMPR117[6] , \A_DOUT_TEMPR118[6] , \A_DOUT_TEMPR0[7] , 
        \A_DOUT_TEMPR1[7] , \A_DOUT_TEMPR2[7] , \A_DOUT_TEMPR3[7] , 
        \A_DOUT_TEMPR4[7] , \A_DOUT_TEMPR5[7] , \A_DOUT_TEMPR6[7] , 
        \A_DOUT_TEMPR7[7] , \A_DOUT_TEMPR8[7] , \A_DOUT_TEMPR9[7] , 
        \A_DOUT_TEMPR10[7] , \A_DOUT_TEMPR11[7] , \A_DOUT_TEMPR12[7] , 
        \A_DOUT_TEMPR13[7] , \A_DOUT_TEMPR14[7] , \A_DOUT_TEMPR15[7] , 
        \A_DOUT_TEMPR16[7] , \A_DOUT_TEMPR17[7] , \A_DOUT_TEMPR18[7] , 
        \A_DOUT_TEMPR19[7] , \A_DOUT_TEMPR20[7] , \A_DOUT_TEMPR21[7] , 
        \A_DOUT_TEMPR22[7] , \A_DOUT_TEMPR23[7] , \A_DOUT_TEMPR24[7] , 
        \A_DOUT_TEMPR25[7] , \A_DOUT_TEMPR26[7] , \A_DOUT_TEMPR27[7] , 
        \A_DOUT_TEMPR28[7] , \A_DOUT_TEMPR29[7] , \A_DOUT_TEMPR30[7] , 
        \A_DOUT_TEMPR31[7] , \A_DOUT_TEMPR32[7] , \A_DOUT_TEMPR33[7] , 
        \A_DOUT_TEMPR34[7] , \A_DOUT_TEMPR35[7] , \A_DOUT_TEMPR36[7] , 
        \A_DOUT_TEMPR37[7] , \A_DOUT_TEMPR38[7] , \A_DOUT_TEMPR39[7] , 
        \A_DOUT_TEMPR40[7] , \A_DOUT_TEMPR41[7] , \A_DOUT_TEMPR42[7] , 
        \A_DOUT_TEMPR43[7] , \A_DOUT_TEMPR44[7] , \A_DOUT_TEMPR45[7] , 
        \A_DOUT_TEMPR46[7] , \A_DOUT_TEMPR47[7] , \A_DOUT_TEMPR48[7] , 
        \A_DOUT_TEMPR49[7] , \A_DOUT_TEMPR50[7] , \A_DOUT_TEMPR51[7] , 
        \A_DOUT_TEMPR52[7] , \A_DOUT_TEMPR53[7] , \A_DOUT_TEMPR54[7] , 
        \A_DOUT_TEMPR55[7] , \A_DOUT_TEMPR56[7] , \A_DOUT_TEMPR57[7] , 
        \A_DOUT_TEMPR58[7] , \A_DOUT_TEMPR59[7] , \A_DOUT_TEMPR60[7] , 
        \A_DOUT_TEMPR61[7] , \A_DOUT_TEMPR62[7] , \A_DOUT_TEMPR63[7] , 
        \A_DOUT_TEMPR64[7] , \A_DOUT_TEMPR65[7] , \A_DOUT_TEMPR66[7] , 
        \A_DOUT_TEMPR67[7] , \A_DOUT_TEMPR68[7] , \A_DOUT_TEMPR69[7] , 
        \A_DOUT_TEMPR70[7] , \A_DOUT_TEMPR71[7] , \A_DOUT_TEMPR72[7] , 
        \A_DOUT_TEMPR73[7] , \A_DOUT_TEMPR74[7] , \A_DOUT_TEMPR75[7] , 
        \A_DOUT_TEMPR76[7] , \A_DOUT_TEMPR77[7] , \A_DOUT_TEMPR78[7] , 
        \A_DOUT_TEMPR79[7] , \A_DOUT_TEMPR80[7] , \A_DOUT_TEMPR81[7] , 
        \A_DOUT_TEMPR82[7] , \A_DOUT_TEMPR83[7] , \A_DOUT_TEMPR84[7] , 
        \A_DOUT_TEMPR85[7] , \A_DOUT_TEMPR86[7] , \A_DOUT_TEMPR87[7] , 
        \A_DOUT_TEMPR88[7] , \A_DOUT_TEMPR89[7] , \A_DOUT_TEMPR90[7] , 
        \A_DOUT_TEMPR91[7] , \A_DOUT_TEMPR92[7] , \A_DOUT_TEMPR93[7] , 
        \A_DOUT_TEMPR94[7] , \A_DOUT_TEMPR95[7] , \A_DOUT_TEMPR96[7] , 
        \A_DOUT_TEMPR97[7] , \A_DOUT_TEMPR98[7] , \A_DOUT_TEMPR99[7] , 
        \A_DOUT_TEMPR100[7] , \A_DOUT_TEMPR101[7] , 
        \A_DOUT_TEMPR102[7] , \A_DOUT_TEMPR103[7] , 
        \A_DOUT_TEMPR104[7] , \A_DOUT_TEMPR105[7] , 
        \A_DOUT_TEMPR106[7] , \A_DOUT_TEMPR107[7] , 
        \A_DOUT_TEMPR108[7] , \A_DOUT_TEMPR109[7] , 
        \A_DOUT_TEMPR110[7] , \A_DOUT_TEMPR111[7] , 
        \A_DOUT_TEMPR112[7] , \A_DOUT_TEMPR113[7] , 
        \A_DOUT_TEMPR114[7] , \A_DOUT_TEMPR115[7] , 
        \A_DOUT_TEMPR116[7] , \A_DOUT_TEMPR117[7] , 
        \A_DOUT_TEMPR118[7] , \A_DOUT_TEMPR0[8] , \A_DOUT_TEMPR1[8] , 
        \A_DOUT_TEMPR2[8] , \A_DOUT_TEMPR3[8] , \A_DOUT_TEMPR4[8] , 
        \A_DOUT_TEMPR5[8] , \A_DOUT_TEMPR6[8] , \A_DOUT_TEMPR7[8] , 
        \A_DOUT_TEMPR8[8] , \A_DOUT_TEMPR9[8] , \A_DOUT_TEMPR10[8] , 
        \A_DOUT_TEMPR11[8] , \A_DOUT_TEMPR12[8] , \A_DOUT_TEMPR13[8] , 
        \A_DOUT_TEMPR14[8] , \A_DOUT_TEMPR15[8] , \A_DOUT_TEMPR16[8] , 
        \A_DOUT_TEMPR17[8] , \A_DOUT_TEMPR18[8] , \A_DOUT_TEMPR19[8] , 
        \A_DOUT_TEMPR20[8] , \A_DOUT_TEMPR21[8] , \A_DOUT_TEMPR22[8] , 
        \A_DOUT_TEMPR23[8] , \A_DOUT_TEMPR24[8] , \A_DOUT_TEMPR25[8] , 
        \A_DOUT_TEMPR26[8] , \A_DOUT_TEMPR27[8] , \A_DOUT_TEMPR28[8] , 
        \A_DOUT_TEMPR29[8] , \A_DOUT_TEMPR30[8] , \A_DOUT_TEMPR31[8] , 
        \A_DOUT_TEMPR32[8] , \A_DOUT_TEMPR33[8] , \A_DOUT_TEMPR34[8] , 
        \A_DOUT_TEMPR35[8] , \A_DOUT_TEMPR36[8] , \A_DOUT_TEMPR37[8] , 
        \A_DOUT_TEMPR38[8] , \A_DOUT_TEMPR39[8] , \A_DOUT_TEMPR40[8] , 
        \A_DOUT_TEMPR41[8] , \A_DOUT_TEMPR42[8] , \A_DOUT_TEMPR43[8] , 
        \A_DOUT_TEMPR44[8] , \A_DOUT_TEMPR45[8] , \A_DOUT_TEMPR46[8] , 
        \A_DOUT_TEMPR47[8] , \A_DOUT_TEMPR48[8] , \A_DOUT_TEMPR49[8] , 
        \A_DOUT_TEMPR50[8] , \A_DOUT_TEMPR51[8] , \A_DOUT_TEMPR52[8] , 
        \A_DOUT_TEMPR53[8] , \A_DOUT_TEMPR54[8] , \A_DOUT_TEMPR55[8] , 
        \A_DOUT_TEMPR56[8] , \A_DOUT_TEMPR57[8] , \A_DOUT_TEMPR58[8] , 
        \A_DOUT_TEMPR59[8] , \A_DOUT_TEMPR60[8] , \A_DOUT_TEMPR61[8] , 
        \A_DOUT_TEMPR62[8] , \A_DOUT_TEMPR63[8] , \A_DOUT_TEMPR64[8] , 
        \A_DOUT_TEMPR65[8] , \A_DOUT_TEMPR66[8] , \A_DOUT_TEMPR67[8] , 
        \A_DOUT_TEMPR68[8] , \A_DOUT_TEMPR69[8] , \A_DOUT_TEMPR70[8] , 
        \A_DOUT_TEMPR71[8] , \A_DOUT_TEMPR72[8] , \A_DOUT_TEMPR73[8] , 
        \A_DOUT_TEMPR74[8] , \A_DOUT_TEMPR75[8] , \A_DOUT_TEMPR76[8] , 
        \A_DOUT_TEMPR77[8] , \A_DOUT_TEMPR78[8] , \A_DOUT_TEMPR79[8] , 
        \A_DOUT_TEMPR80[8] , \A_DOUT_TEMPR81[8] , \A_DOUT_TEMPR82[8] , 
        \A_DOUT_TEMPR83[8] , \A_DOUT_TEMPR84[8] , \A_DOUT_TEMPR85[8] , 
        \A_DOUT_TEMPR86[8] , \A_DOUT_TEMPR87[8] , \A_DOUT_TEMPR88[8] , 
        \A_DOUT_TEMPR89[8] , \A_DOUT_TEMPR90[8] , \A_DOUT_TEMPR91[8] , 
        \A_DOUT_TEMPR92[8] , \A_DOUT_TEMPR93[8] , \A_DOUT_TEMPR94[8] , 
        \A_DOUT_TEMPR95[8] , \A_DOUT_TEMPR96[8] , \A_DOUT_TEMPR97[8] , 
        \A_DOUT_TEMPR98[8] , \A_DOUT_TEMPR99[8] , \A_DOUT_TEMPR100[8] , 
        \A_DOUT_TEMPR101[8] , \A_DOUT_TEMPR102[8] , 
        \A_DOUT_TEMPR103[8] , \A_DOUT_TEMPR104[8] , 
        \A_DOUT_TEMPR105[8] , \A_DOUT_TEMPR106[8] , 
        \A_DOUT_TEMPR107[8] , \A_DOUT_TEMPR108[8] , 
        \A_DOUT_TEMPR109[8] , \A_DOUT_TEMPR110[8] , 
        \A_DOUT_TEMPR111[8] , \A_DOUT_TEMPR112[8] , 
        \A_DOUT_TEMPR113[8] , \A_DOUT_TEMPR114[8] , 
        \A_DOUT_TEMPR115[8] , \A_DOUT_TEMPR116[8] , 
        \A_DOUT_TEMPR117[8] , \A_DOUT_TEMPR118[8] , \A_DOUT_TEMPR0[9] , 
        \A_DOUT_TEMPR1[9] , \A_DOUT_TEMPR2[9] , \A_DOUT_TEMPR3[9] , 
        \A_DOUT_TEMPR4[9] , \A_DOUT_TEMPR5[9] , \A_DOUT_TEMPR6[9] , 
        \A_DOUT_TEMPR7[9] , \A_DOUT_TEMPR8[9] , \A_DOUT_TEMPR9[9] , 
        \A_DOUT_TEMPR10[9] , \A_DOUT_TEMPR11[9] , \A_DOUT_TEMPR12[9] , 
        \A_DOUT_TEMPR13[9] , \A_DOUT_TEMPR14[9] , \A_DOUT_TEMPR15[9] , 
        \A_DOUT_TEMPR16[9] , \A_DOUT_TEMPR17[9] , \A_DOUT_TEMPR18[9] , 
        \A_DOUT_TEMPR19[9] , \A_DOUT_TEMPR20[9] , \A_DOUT_TEMPR21[9] , 
        \A_DOUT_TEMPR22[9] , \A_DOUT_TEMPR23[9] , \A_DOUT_TEMPR24[9] , 
        \A_DOUT_TEMPR25[9] , \A_DOUT_TEMPR26[9] , \A_DOUT_TEMPR27[9] , 
        \A_DOUT_TEMPR28[9] , \A_DOUT_TEMPR29[9] , \A_DOUT_TEMPR30[9] , 
        \A_DOUT_TEMPR31[9] , \A_DOUT_TEMPR32[9] , \A_DOUT_TEMPR33[9] , 
        \A_DOUT_TEMPR34[9] , \A_DOUT_TEMPR35[9] , \A_DOUT_TEMPR36[9] , 
        \A_DOUT_TEMPR37[9] , \A_DOUT_TEMPR38[9] , \A_DOUT_TEMPR39[9] , 
        \A_DOUT_TEMPR40[9] , \A_DOUT_TEMPR41[9] , \A_DOUT_TEMPR42[9] , 
        \A_DOUT_TEMPR43[9] , \A_DOUT_TEMPR44[9] , \A_DOUT_TEMPR45[9] , 
        \A_DOUT_TEMPR46[9] , \A_DOUT_TEMPR47[9] , \A_DOUT_TEMPR48[9] , 
        \A_DOUT_TEMPR49[9] , \A_DOUT_TEMPR50[9] , \A_DOUT_TEMPR51[9] , 
        \A_DOUT_TEMPR52[9] , \A_DOUT_TEMPR53[9] , \A_DOUT_TEMPR54[9] , 
        \A_DOUT_TEMPR55[9] , \A_DOUT_TEMPR56[9] , \A_DOUT_TEMPR57[9] , 
        \A_DOUT_TEMPR58[9] , \A_DOUT_TEMPR59[9] , \A_DOUT_TEMPR60[9] , 
        \A_DOUT_TEMPR61[9] , \A_DOUT_TEMPR62[9] , \A_DOUT_TEMPR63[9] , 
        \A_DOUT_TEMPR64[9] , \A_DOUT_TEMPR65[9] , \A_DOUT_TEMPR66[9] , 
        \A_DOUT_TEMPR67[9] , \A_DOUT_TEMPR68[9] , \A_DOUT_TEMPR69[9] , 
        \A_DOUT_TEMPR70[9] , \A_DOUT_TEMPR71[9] , \A_DOUT_TEMPR72[9] , 
        \A_DOUT_TEMPR73[9] , \A_DOUT_TEMPR74[9] , \A_DOUT_TEMPR75[9] , 
        \A_DOUT_TEMPR76[9] , \A_DOUT_TEMPR77[9] , \A_DOUT_TEMPR78[9] , 
        \A_DOUT_TEMPR79[9] , \A_DOUT_TEMPR80[9] , \A_DOUT_TEMPR81[9] , 
        \A_DOUT_TEMPR82[9] , \A_DOUT_TEMPR83[9] , \A_DOUT_TEMPR84[9] , 
        \A_DOUT_TEMPR85[9] , \A_DOUT_TEMPR86[9] , \A_DOUT_TEMPR87[9] , 
        \A_DOUT_TEMPR88[9] , \A_DOUT_TEMPR89[9] , \A_DOUT_TEMPR90[9] , 
        \A_DOUT_TEMPR91[9] , \A_DOUT_TEMPR92[9] , \A_DOUT_TEMPR93[9] , 
        \A_DOUT_TEMPR94[9] , \A_DOUT_TEMPR95[9] , \A_DOUT_TEMPR96[9] , 
        \A_DOUT_TEMPR97[9] , \A_DOUT_TEMPR98[9] , \A_DOUT_TEMPR99[9] , 
        \A_DOUT_TEMPR100[9] , \A_DOUT_TEMPR101[9] , 
        \A_DOUT_TEMPR102[9] , \A_DOUT_TEMPR103[9] , 
        \A_DOUT_TEMPR104[9] , \A_DOUT_TEMPR105[9] , 
        \A_DOUT_TEMPR106[9] , \A_DOUT_TEMPR107[9] , 
        \A_DOUT_TEMPR108[9] , \A_DOUT_TEMPR109[9] , 
        \A_DOUT_TEMPR110[9] , \A_DOUT_TEMPR111[9] , 
        \A_DOUT_TEMPR112[9] , \A_DOUT_TEMPR113[9] , 
        \A_DOUT_TEMPR114[9] , \A_DOUT_TEMPR115[9] , 
        \A_DOUT_TEMPR116[9] , \A_DOUT_TEMPR117[9] , 
        \A_DOUT_TEMPR118[9] , \A_DOUT_TEMPR0[10] , \A_DOUT_TEMPR1[10] , 
        \A_DOUT_TEMPR2[10] , \A_DOUT_TEMPR3[10] , \A_DOUT_TEMPR4[10] , 
        \A_DOUT_TEMPR5[10] , \A_DOUT_TEMPR6[10] , \A_DOUT_TEMPR7[10] , 
        \A_DOUT_TEMPR8[10] , \A_DOUT_TEMPR9[10] , \A_DOUT_TEMPR10[10] , 
        \A_DOUT_TEMPR11[10] , \A_DOUT_TEMPR12[10] , 
        \A_DOUT_TEMPR13[10] , \A_DOUT_TEMPR14[10] , 
        \A_DOUT_TEMPR15[10] , \A_DOUT_TEMPR16[10] , 
        \A_DOUT_TEMPR17[10] , \A_DOUT_TEMPR18[10] , 
        \A_DOUT_TEMPR19[10] , \A_DOUT_TEMPR20[10] , 
        \A_DOUT_TEMPR21[10] , \A_DOUT_TEMPR22[10] , 
        \A_DOUT_TEMPR23[10] , \A_DOUT_TEMPR24[10] , 
        \A_DOUT_TEMPR25[10] , \A_DOUT_TEMPR26[10] , 
        \A_DOUT_TEMPR27[10] , \A_DOUT_TEMPR28[10] , 
        \A_DOUT_TEMPR29[10] , \A_DOUT_TEMPR30[10] , 
        \A_DOUT_TEMPR31[10] , \A_DOUT_TEMPR32[10] , 
        \A_DOUT_TEMPR33[10] , \A_DOUT_TEMPR34[10] , 
        \A_DOUT_TEMPR35[10] , \A_DOUT_TEMPR36[10] , 
        \A_DOUT_TEMPR37[10] , \A_DOUT_TEMPR38[10] , 
        \A_DOUT_TEMPR39[10] , \A_DOUT_TEMPR40[10] , 
        \A_DOUT_TEMPR41[10] , \A_DOUT_TEMPR42[10] , 
        \A_DOUT_TEMPR43[10] , \A_DOUT_TEMPR44[10] , 
        \A_DOUT_TEMPR45[10] , \A_DOUT_TEMPR46[10] , 
        \A_DOUT_TEMPR47[10] , \A_DOUT_TEMPR48[10] , 
        \A_DOUT_TEMPR49[10] , \A_DOUT_TEMPR50[10] , 
        \A_DOUT_TEMPR51[10] , \A_DOUT_TEMPR52[10] , 
        \A_DOUT_TEMPR53[10] , \A_DOUT_TEMPR54[10] , 
        \A_DOUT_TEMPR55[10] , \A_DOUT_TEMPR56[10] , 
        \A_DOUT_TEMPR57[10] , \A_DOUT_TEMPR58[10] , 
        \A_DOUT_TEMPR59[10] , \A_DOUT_TEMPR60[10] , 
        \A_DOUT_TEMPR61[10] , \A_DOUT_TEMPR62[10] , 
        \A_DOUT_TEMPR63[10] , \A_DOUT_TEMPR64[10] , 
        \A_DOUT_TEMPR65[10] , \A_DOUT_TEMPR66[10] , 
        \A_DOUT_TEMPR67[10] , \A_DOUT_TEMPR68[10] , 
        \A_DOUT_TEMPR69[10] , \A_DOUT_TEMPR70[10] , 
        \A_DOUT_TEMPR71[10] , \A_DOUT_TEMPR72[10] , 
        \A_DOUT_TEMPR73[10] , \A_DOUT_TEMPR74[10] , 
        \A_DOUT_TEMPR75[10] , \A_DOUT_TEMPR76[10] , 
        \A_DOUT_TEMPR77[10] , \A_DOUT_TEMPR78[10] , 
        \A_DOUT_TEMPR79[10] , \A_DOUT_TEMPR80[10] , 
        \A_DOUT_TEMPR81[10] , \A_DOUT_TEMPR82[10] , 
        \A_DOUT_TEMPR83[10] , \A_DOUT_TEMPR84[10] , 
        \A_DOUT_TEMPR85[10] , \A_DOUT_TEMPR86[10] , 
        \A_DOUT_TEMPR87[10] , \A_DOUT_TEMPR88[10] , 
        \A_DOUT_TEMPR89[10] , \A_DOUT_TEMPR90[10] , 
        \A_DOUT_TEMPR91[10] , \A_DOUT_TEMPR92[10] , 
        \A_DOUT_TEMPR93[10] , \A_DOUT_TEMPR94[10] , 
        \A_DOUT_TEMPR95[10] , \A_DOUT_TEMPR96[10] , 
        \A_DOUT_TEMPR97[10] , \A_DOUT_TEMPR98[10] , 
        \A_DOUT_TEMPR99[10] , \A_DOUT_TEMPR100[10] , 
        \A_DOUT_TEMPR101[10] , \A_DOUT_TEMPR102[10] , 
        \A_DOUT_TEMPR103[10] , \A_DOUT_TEMPR104[10] , 
        \A_DOUT_TEMPR105[10] , \A_DOUT_TEMPR106[10] , 
        \A_DOUT_TEMPR107[10] , \A_DOUT_TEMPR108[10] , 
        \A_DOUT_TEMPR109[10] , \A_DOUT_TEMPR110[10] , 
        \A_DOUT_TEMPR111[10] , \A_DOUT_TEMPR112[10] , 
        \A_DOUT_TEMPR113[10] , \A_DOUT_TEMPR114[10] , 
        \A_DOUT_TEMPR115[10] , \A_DOUT_TEMPR116[10] , 
        \A_DOUT_TEMPR117[10] , \A_DOUT_TEMPR118[10] , 
        \A_DOUT_TEMPR0[11] , \A_DOUT_TEMPR1[11] , \A_DOUT_TEMPR2[11] , 
        \A_DOUT_TEMPR3[11] , \A_DOUT_TEMPR4[11] , \A_DOUT_TEMPR5[11] , 
        \A_DOUT_TEMPR6[11] , \A_DOUT_TEMPR7[11] , \A_DOUT_TEMPR8[11] , 
        \A_DOUT_TEMPR9[11] , \A_DOUT_TEMPR10[11] , 
        \A_DOUT_TEMPR11[11] , \A_DOUT_TEMPR12[11] , 
        \A_DOUT_TEMPR13[11] , \A_DOUT_TEMPR14[11] , 
        \A_DOUT_TEMPR15[11] , \A_DOUT_TEMPR16[11] , 
        \A_DOUT_TEMPR17[11] , \A_DOUT_TEMPR18[11] , 
        \A_DOUT_TEMPR19[11] , \A_DOUT_TEMPR20[11] , 
        \A_DOUT_TEMPR21[11] , \A_DOUT_TEMPR22[11] , 
        \A_DOUT_TEMPR23[11] , \A_DOUT_TEMPR24[11] , 
        \A_DOUT_TEMPR25[11] , \A_DOUT_TEMPR26[11] , 
        \A_DOUT_TEMPR27[11] , \A_DOUT_TEMPR28[11] , 
        \A_DOUT_TEMPR29[11] , \A_DOUT_TEMPR30[11] , 
        \A_DOUT_TEMPR31[11] , \A_DOUT_TEMPR32[11] , 
        \A_DOUT_TEMPR33[11] , \A_DOUT_TEMPR34[11] , 
        \A_DOUT_TEMPR35[11] , \A_DOUT_TEMPR36[11] , 
        \A_DOUT_TEMPR37[11] , \A_DOUT_TEMPR38[11] , 
        \A_DOUT_TEMPR39[11] , \A_DOUT_TEMPR40[11] , 
        \A_DOUT_TEMPR41[11] , \A_DOUT_TEMPR42[11] , 
        \A_DOUT_TEMPR43[11] , \A_DOUT_TEMPR44[11] , 
        \A_DOUT_TEMPR45[11] , \A_DOUT_TEMPR46[11] , 
        \A_DOUT_TEMPR47[11] , \A_DOUT_TEMPR48[11] , 
        \A_DOUT_TEMPR49[11] , \A_DOUT_TEMPR50[11] , 
        \A_DOUT_TEMPR51[11] , \A_DOUT_TEMPR52[11] , 
        \A_DOUT_TEMPR53[11] , \A_DOUT_TEMPR54[11] , 
        \A_DOUT_TEMPR55[11] , \A_DOUT_TEMPR56[11] , 
        \A_DOUT_TEMPR57[11] , \A_DOUT_TEMPR58[11] , 
        \A_DOUT_TEMPR59[11] , \A_DOUT_TEMPR60[11] , 
        \A_DOUT_TEMPR61[11] , \A_DOUT_TEMPR62[11] , 
        \A_DOUT_TEMPR63[11] , \A_DOUT_TEMPR64[11] , 
        \A_DOUT_TEMPR65[11] , \A_DOUT_TEMPR66[11] , 
        \A_DOUT_TEMPR67[11] , \A_DOUT_TEMPR68[11] , 
        \A_DOUT_TEMPR69[11] , \A_DOUT_TEMPR70[11] , 
        \A_DOUT_TEMPR71[11] , \A_DOUT_TEMPR72[11] , 
        \A_DOUT_TEMPR73[11] , \A_DOUT_TEMPR74[11] , 
        \A_DOUT_TEMPR75[11] , \A_DOUT_TEMPR76[11] , 
        \A_DOUT_TEMPR77[11] , \A_DOUT_TEMPR78[11] , 
        \A_DOUT_TEMPR79[11] , \A_DOUT_TEMPR80[11] , 
        \A_DOUT_TEMPR81[11] , \A_DOUT_TEMPR82[11] , 
        \A_DOUT_TEMPR83[11] , \A_DOUT_TEMPR84[11] , 
        \A_DOUT_TEMPR85[11] , \A_DOUT_TEMPR86[11] , 
        \A_DOUT_TEMPR87[11] , \A_DOUT_TEMPR88[11] , 
        \A_DOUT_TEMPR89[11] , \A_DOUT_TEMPR90[11] , 
        \A_DOUT_TEMPR91[11] , \A_DOUT_TEMPR92[11] , 
        \A_DOUT_TEMPR93[11] , \A_DOUT_TEMPR94[11] , 
        \A_DOUT_TEMPR95[11] , \A_DOUT_TEMPR96[11] , 
        \A_DOUT_TEMPR97[11] , \A_DOUT_TEMPR98[11] , 
        \A_DOUT_TEMPR99[11] , \A_DOUT_TEMPR100[11] , 
        \A_DOUT_TEMPR101[11] , \A_DOUT_TEMPR102[11] , 
        \A_DOUT_TEMPR103[11] , \A_DOUT_TEMPR104[11] , 
        \A_DOUT_TEMPR105[11] , \A_DOUT_TEMPR106[11] , 
        \A_DOUT_TEMPR107[11] , \A_DOUT_TEMPR108[11] , 
        \A_DOUT_TEMPR109[11] , \A_DOUT_TEMPR110[11] , 
        \A_DOUT_TEMPR111[11] , \A_DOUT_TEMPR112[11] , 
        \A_DOUT_TEMPR113[11] , \A_DOUT_TEMPR114[11] , 
        \A_DOUT_TEMPR115[11] , \A_DOUT_TEMPR116[11] , 
        \A_DOUT_TEMPR117[11] , \A_DOUT_TEMPR118[11] , 
        \A_DOUT_TEMPR0[12] , \A_DOUT_TEMPR1[12] , \A_DOUT_TEMPR2[12] , 
        \A_DOUT_TEMPR3[12] , \A_DOUT_TEMPR4[12] , \A_DOUT_TEMPR5[12] , 
        \A_DOUT_TEMPR6[12] , \A_DOUT_TEMPR7[12] , \A_DOUT_TEMPR8[12] , 
        \A_DOUT_TEMPR9[12] , \A_DOUT_TEMPR10[12] , 
        \A_DOUT_TEMPR11[12] , \A_DOUT_TEMPR12[12] , 
        \A_DOUT_TEMPR13[12] , \A_DOUT_TEMPR14[12] , 
        \A_DOUT_TEMPR15[12] , \A_DOUT_TEMPR16[12] , 
        \A_DOUT_TEMPR17[12] , \A_DOUT_TEMPR18[12] , 
        \A_DOUT_TEMPR19[12] , \A_DOUT_TEMPR20[12] , 
        \A_DOUT_TEMPR21[12] , \A_DOUT_TEMPR22[12] , 
        \A_DOUT_TEMPR23[12] , \A_DOUT_TEMPR24[12] , 
        \A_DOUT_TEMPR25[12] , \A_DOUT_TEMPR26[12] , 
        \A_DOUT_TEMPR27[12] , \A_DOUT_TEMPR28[12] , 
        \A_DOUT_TEMPR29[12] , \A_DOUT_TEMPR30[12] , 
        \A_DOUT_TEMPR31[12] , \A_DOUT_TEMPR32[12] , 
        \A_DOUT_TEMPR33[12] , \A_DOUT_TEMPR34[12] , 
        \A_DOUT_TEMPR35[12] , \A_DOUT_TEMPR36[12] , 
        \A_DOUT_TEMPR37[12] , \A_DOUT_TEMPR38[12] , 
        \A_DOUT_TEMPR39[12] , \A_DOUT_TEMPR40[12] , 
        \A_DOUT_TEMPR41[12] , \A_DOUT_TEMPR42[12] , 
        \A_DOUT_TEMPR43[12] , \A_DOUT_TEMPR44[12] , 
        \A_DOUT_TEMPR45[12] , \A_DOUT_TEMPR46[12] , 
        \A_DOUT_TEMPR47[12] , \A_DOUT_TEMPR48[12] , 
        \A_DOUT_TEMPR49[12] , \A_DOUT_TEMPR50[12] , 
        \A_DOUT_TEMPR51[12] , \A_DOUT_TEMPR52[12] , 
        \A_DOUT_TEMPR53[12] , \A_DOUT_TEMPR54[12] , 
        \A_DOUT_TEMPR55[12] , \A_DOUT_TEMPR56[12] , 
        \A_DOUT_TEMPR57[12] , \A_DOUT_TEMPR58[12] , 
        \A_DOUT_TEMPR59[12] , \A_DOUT_TEMPR60[12] , 
        \A_DOUT_TEMPR61[12] , \A_DOUT_TEMPR62[12] , 
        \A_DOUT_TEMPR63[12] , \A_DOUT_TEMPR64[12] , 
        \A_DOUT_TEMPR65[12] , \A_DOUT_TEMPR66[12] , 
        \A_DOUT_TEMPR67[12] , \A_DOUT_TEMPR68[12] , 
        \A_DOUT_TEMPR69[12] , \A_DOUT_TEMPR70[12] , 
        \A_DOUT_TEMPR71[12] , \A_DOUT_TEMPR72[12] , 
        \A_DOUT_TEMPR73[12] , \A_DOUT_TEMPR74[12] , 
        \A_DOUT_TEMPR75[12] , \A_DOUT_TEMPR76[12] , 
        \A_DOUT_TEMPR77[12] , \A_DOUT_TEMPR78[12] , 
        \A_DOUT_TEMPR79[12] , \A_DOUT_TEMPR80[12] , 
        \A_DOUT_TEMPR81[12] , \A_DOUT_TEMPR82[12] , 
        \A_DOUT_TEMPR83[12] , \A_DOUT_TEMPR84[12] , 
        \A_DOUT_TEMPR85[12] , \A_DOUT_TEMPR86[12] , 
        \A_DOUT_TEMPR87[12] , \A_DOUT_TEMPR88[12] , 
        \A_DOUT_TEMPR89[12] , \A_DOUT_TEMPR90[12] , 
        \A_DOUT_TEMPR91[12] , \A_DOUT_TEMPR92[12] , 
        \A_DOUT_TEMPR93[12] , \A_DOUT_TEMPR94[12] , 
        \A_DOUT_TEMPR95[12] , \A_DOUT_TEMPR96[12] , 
        \A_DOUT_TEMPR97[12] , \A_DOUT_TEMPR98[12] , 
        \A_DOUT_TEMPR99[12] , \A_DOUT_TEMPR100[12] , 
        \A_DOUT_TEMPR101[12] , \A_DOUT_TEMPR102[12] , 
        \A_DOUT_TEMPR103[12] , \A_DOUT_TEMPR104[12] , 
        \A_DOUT_TEMPR105[12] , \A_DOUT_TEMPR106[12] , 
        \A_DOUT_TEMPR107[12] , \A_DOUT_TEMPR108[12] , 
        \A_DOUT_TEMPR109[12] , \A_DOUT_TEMPR110[12] , 
        \A_DOUT_TEMPR111[12] , \A_DOUT_TEMPR112[12] , 
        \A_DOUT_TEMPR113[12] , \A_DOUT_TEMPR114[12] , 
        \A_DOUT_TEMPR115[12] , \A_DOUT_TEMPR116[12] , 
        \A_DOUT_TEMPR117[12] , \A_DOUT_TEMPR118[12] , 
        \A_DOUT_TEMPR0[13] , \A_DOUT_TEMPR1[13] , \A_DOUT_TEMPR2[13] , 
        \A_DOUT_TEMPR3[13] , \A_DOUT_TEMPR4[13] , \A_DOUT_TEMPR5[13] , 
        \A_DOUT_TEMPR6[13] , \A_DOUT_TEMPR7[13] , \A_DOUT_TEMPR8[13] , 
        \A_DOUT_TEMPR9[13] , \A_DOUT_TEMPR10[13] , 
        \A_DOUT_TEMPR11[13] , \A_DOUT_TEMPR12[13] , 
        \A_DOUT_TEMPR13[13] , \A_DOUT_TEMPR14[13] , 
        \A_DOUT_TEMPR15[13] , \A_DOUT_TEMPR16[13] , 
        \A_DOUT_TEMPR17[13] , \A_DOUT_TEMPR18[13] , 
        \A_DOUT_TEMPR19[13] , \A_DOUT_TEMPR20[13] , 
        \A_DOUT_TEMPR21[13] , \A_DOUT_TEMPR22[13] , 
        \A_DOUT_TEMPR23[13] , \A_DOUT_TEMPR24[13] , 
        \A_DOUT_TEMPR25[13] , \A_DOUT_TEMPR26[13] , 
        \A_DOUT_TEMPR27[13] , \A_DOUT_TEMPR28[13] , 
        \A_DOUT_TEMPR29[13] , \A_DOUT_TEMPR30[13] , 
        \A_DOUT_TEMPR31[13] , \A_DOUT_TEMPR32[13] , 
        \A_DOUT_TEMPR33[13] , \A_DOUT_TEMPR34[13] , 
        \A_DOUT_TEMPR35[13] , \A_DOUT_TEMPR36[13] , 
        \A_DOUT_TEMPR37[13] , \A_DOUT_TEMPR38[13] , 
        \A_DOUT_TEMPR39[13] , \A_DOUT_TEMPR40[13] , 
        \A_DOUT_TEMPR41[13] , \A_DOUT_TEMPR42[13] , 
        \A_DOUT_TEMPR43[13] , \A_DOUT_TEMPR44[13] , 
        \A_DOUT_TEMPR45[13] , \A_DOUT_TEMPR46[13] , 
        \A_DOUT_TEMPR47[13] , \A_DOUT_TEMPR48[13] , 
        \A_DOUT_TEMPR49[13] , \A_DOUT_TEMPR50[13] , 
        \A_DOUT_TEMPR51[13] , \A_DOUT_TEMPR52[13] , 
        \A_DOUT_TEMPR53[13] , \A_DOUT_TEMPR54[13] , 
        \A_DOUT_TEMPR55[13] , \A_DOUT_TEMPR56[13] , 
        \A_DOUT_TEMPR57[13] , \A_DOUT_TEMPR58[13] , 
        \A_DOUT_TEMPR59[13] , \A_DOUT_TEMPR60[13] , 
        \A_DOUT_TEMPR61[13] , \A_DOUT_TEMPR62[13] , 
        \A_DOUT_TEMPR63[13] , \A_DOUT_TEMPR64[13] , 
        \A_DOUT_TEMPR65[13] , \A_DOUT_TEMPR66[13] , 
        \A_DOUT_TEMPR67[13] , \A_DOUT_TEMPR68[13] , 
        \A_DOUT_TEMPR69[13] , \A_DOUT_TEMPR70[13] , 
        \A_DOUT_TEMPR71[13] , \A_DOUT_TEMPR72[13] , 
        \A_DOUT_TEMPR73[13] , \A_DOUT_TEMPR74[13] , 
        \A_DOUT_TEMPR75[13] , \A_DOUT_TEMPR76[13] , 
        \A_DOUT_TEMPR77[13] , \A_DOUT_TEMPR78[13] , 
        \A_DOUT_TEMPR79[13] , \A_DOUT_TEMPR80[13] , 
        \A_DOUT_TEMPR81[13] , \A_DOUT_TEMPR82[13] , 
        \A_DOUT_TEMPR83[13] , \A_DOUT_TEMPR84[13] , 
        \A_DOUT_TEMPR85[13] , \A_DOUT_TEMPR86[13] , 
        \A_DOUT_TEMPR87[13] , \A_DOUT_TEMPR88[13] , 
        \A_DOUT_TEMPR89[13] , \A_DOUT_TEMPR90[13] , 
        \A_DOUT_TEMPR91[13] , \A_DOUT_TEMPR92[13] , 
        \A_DOUT_TEMPR93[13] , \A_DOUT_TEMPR94[13] , 
        \A_DOUT_TEMPR95[13] , \A_DOUT_TEMPR96[13] , 
        \A_DOUT_TEMPR97[13] , \A_DOUT_TEMPR98[13] , 
        \A_DOUT_TEMPR99[13] , \A_DOUT_TEMPR100[13] , 
        \A_DOUT_TEMPR101[13] , \A_DOUT_TEMPR102[13] , 
        \A_DOUT_TEMPR103[13] , \A_DOUT_TEMPR104[13] , 
        \A_DOUT_TEMPR105[13] , \A_DOUT_TEMPR106[13] , 
        \A_DOUT_TEMPR107[13] , \A_DOUT_TEMPR108[13] , 
        \A_DOUT_TEMPR109[13] , \A_DOUT_TEMPR110[13] , 
        \A_DOUT_TEMPR111[13] , \A_DOUT_TEMPR112[13] , 
        \A_DOUT_TEMPR113[13] , \A_DOUT_TEMPR114[13] , 
        \A_DOUT_TEMPR115[13] , \A_DOUT_TEMPR116[13] , 
        \A_DOUT_TEMPR117[13] , \A_DOUT_TEMPR118[13] , 
        \A_DOUT_TEMPR0[14] , \A_DOUT_TEMPR1[14] , \A_DOUT_TEMPR2[14] , 
        \A_DOUT_TEMPR3[14] , \A_DOUT_TEMPR4[14] , \A_DOUT_TEMPR5[14] , 
        \A_DOUT_TEMPR6[14] , \A_DOUT_TEMPR7[14] , \A_DOUT_TEMPR8[14] , 
        \A_DOUT_TEMPR9[14] , \A_DOUT_TEMPR10[14] , 
        \A_DOUT_TEMPR11[14] , \A_DOUT_TEMPR12[14] , 
        \A_DOUT_TEMPR13[14] , \A_DOUT_TEMPR14[14] , 
        \A_DOUT_TEMPR15[14] , \A_DOUT_TEMPR16[14] , 
        \A_DOUT_TEMPR17[14] , \A_DOUT_TEMPR18[14] , 
        \A_DOUT_TEMPR19[14] , \A_DOUT_TEMPR20[14] , 
        \A_DOUT_TEMPR21[14] , \A_DOUT_TEMPR22[14] , 
        \A_DOUT_TEMPR23[14] , \A_DOUT_TEMPR24[14] , 
        \A_DOUT_TEMPR25[14] , \A_DOUT_TEMPR26[14] , 
        \A_DOUT_TEMPR27[14] , \A_DOUT_TEMPR28[14] , 
        \A_DOUT_TEMPR29[14] , \A_DOUT_TEMPR30[14] , 
        \A_DOUT_TEMPR31[14] , \A_DOUT_TEMPR32[14] , 
        \A_DOUT_TEMPR33[14] , \A_DOUT_TEMPR34[14] , 
        \A_DOUT_TEMPR35[14] , \A_DOUT_TEMPR36[14] , 
        \A_DOUT_TEMPR37[14] , \A_DOUT_TEMPR38[14] , 
        \A_DOUT_TEMPR39[14] , \A_DOUT_TEMPR40[14] , 
        \A_DOUT_TEMPR41[14] , \A_DOUT_TEMPR42[14] , 
        \A_DOUT_TEMPR43[14] , \A_DOUT_TEMPR44[14] , 
        \A_DOUT_TEMPR45[14] , \A_DOUT_TEMPR46[14] , 
        \A_DOUT_TEMPR47[14] , \A_DOUT_TEMPR48[14] , 
        \A_DOUT_TEMPR49[14] , \A_DOUT_TEMPR50[14] , 
        \A_DOUT_TEMPR51[14] , \A_DOUT_TEMPR52[14] , 
        \A_DOUT_TEMPR53[14] , \A_DOUT_TEMPR54[14] , 
        \A_DOUT_TEMPR55[14] , \A_DOUT_TEMPR56[14] , 
        \A_DOUT_TEMPR57[14] , \A_DOUT_TEMPR58[14] , 
        \A_DOUT_TEMPR59[14] , \A_DOUT_TEMPR60[14] , 
        \A_DOUT_TEMPR61[14] , \A_DOUT_TEMPR62[14] , 
        \A_DOUT_TEMPR63[14] , \A_DOUT_TEMPR64[14] , 
        \A_DOUT_TEMPR65[14] , \A_DOUT_TEMPR66[14] , 
        \A_DOUT_TEMPR67[14] , \A_DOUT_TEMPR68[14] , 
        \A_DOUT_TEMPR69[14] , \A_DOUT_TEMPR70[14] , 
        \A_DOUT_TEMPR71[14] , \A_DOUT_TEMPR72[14] , 
        \A_DOUT_TEMPR73[14] , \A_DOUT_TEMPR74[14] , 
        \A_DOUT_TEMPR75[14] , \A_DOUT_TEMPR76[14] , 
        \A_DOUT_TEMPR77[14] , \A_DOUT_TEMPR78[14] , 
        \A_DOUT_TEMPR79[14] , \A_DOUT_TEMPR80[14] , 
        \A_DOUT_TEMPR81[14] , \A_DOUT_TEMPR82[14] , 
        \A_DOUT_TEMPR83[14] , \A_DOUT_TEMPR84[14] , 
        \A_DOUT_TEMPR85[14] , \A_DOUT_TEMPR86[14] , 
        \A_DOUT_TEMPR87[14] , \A_DOUT_TEMPR88[14] , 
        \A_DOUT_TEMPR89[14] , \A_DOUT_TEMPR90[14] , 
        \A_DOUT_TEMPR91[14] , \A_DOUT_TEMPR92[14] , 
        \A_DOUT_TEMPR93[14] , \A_DOUT_TEMPR94[14] , 
        \A_DOUT_TEMPR95[14] , \A_DOUT_TEMPR96[14] , 
        \A_DOUT_TEMPR97[14] , \A_DOUT_TEMPR98[14] , 
        \A_DOUT_TEMPR99[14] , \A_DOUT_TEMPR100[14] , 
        \A_DOUT_TEMPR101[14] , \A_DOUT_TEMPR102[14] , 
        \A_DOUT_TEMPR103[14] , \A_DOUT_TEMPR104[14] , 
        \A_DOUT_TEMPR105[14] , \A_DOUT_TEMPR106[14] , 
        \A_DOUT_TEMPR107[14] , \A_DOUT_TEMPR108[14] , 
        \A_DOUT_TEMPR109[14] , \A_DOUT_TEMPR110[14] , 
        \A_DOUT_TEMPR111[14] , \A_DOUT_TEMPR112[14] , 
        \A_DOUT_TEMPR113[14] , \A_DOUT_TEMPR114[14] , 
        \A_DOUT_TEMPR115[14] , \A_DOUT_TEMPR116[14] , 
        \A_DOUT_TEMPR117[14] , \A_DOUT_TEMPR118[14] , 
        \A_DOUT_TEMPR0[15] , \A_DOUT_TEMPR1[15] , \A_DOUT_TEMPR2[15] , 
        \A_DOUT_TEMPR3[15] , \A_DOUT_TEMPR4[15] , \A_DOUT_TEMPR5[15] , 
        \A_DOUT_TEMPR6[15] , \A_DOUT_TEMPR7[15] , \A_DOUT_TEMPR8[15] , 
        \A_DOUT_TEMPR9[15] , \A_DOUT_TEMPR10[15] , 
        \A_DOUT_TEMPR11[15] , \A_DOUT_TEMPR12[15] , 
        \A_DOUT_TEMPR13[15] , \A_DOUT_TEMPR14[15] , 
        \A_DOUT_TEMPR15[15] , \A_DOUT_TEMPR16[15] , 
        \A_DOUT_TEMPR17[15] , \A_DOUT_TEMPR18[15] , 
        \A_DOUT_TEMPR19[15] , \A_DOUT_TEMPR20[15] , 
        \A_DOUT_TEMPR21[15] , \A_DOUT_TEMPR22[15] , 
        \A_DOUT_TEMPR23[15] , \A_DOUT_TEMPR24[15] , 
        \A_DOUT_TEMPR25[15] , \A_DOUT_TEMPR26[15] , 
        \A_DOUT_TEMPR27[15] , \A_DOUT_TEMPR28[15] , 
        \A_DOUT_TEMPR29[15] , \A_DOUT_TEMPR30[15] , 
        \A_DOUT_TEMPR31[15] , \A_DOUT_TEMPR32[15] , 
        \A_DOUT_TEMPR33[15] , \A_DOUT_TEMPR34[15] , 
        \A_DOUT_TEMPR35[15] , \A_DOUT_TEMPR36[15] , 
        \A_DOUT_TEMPR37[15] , \A_DOUT_TEMPR38[15] , 
        \A_DOUT_TEMPR39[15] , \A_DOUT_TEMPR40[15] , 
        \A_DOUT_TEMPR41[15] , \A_DOUT_TEMPR42[15] , 
        \A_DOUT_TEMPR43[15] , \A_DOUT_TEMPR44[15] , 
        \A_DOUT_TEMPR45[15] , \A_DOUT_TEMPR46[15] , 
        \A_DOUT_TEMPR47[15] , \A_DOUT_TEMPR48[15] , 
        \A_DOUT_TEMPR49[15] , \A_DOUT_TEMPR50[15] , 
        \A_DOUT_TEMPR51[15] , \A_DOUT_TEMPR52[15] , 
        \A_DOUT_TEMPR53[15] , \A_DOUT_TEMPR54[15] , 
        \A_DOUT_TEMPR55[15] , \A_DOUT_TEMPR56[15] , 
        \A_DOUT_TEMPR57[15] , \A_DOUT_TEMPR58[15] , 
        \A_DOUT_TEMPR59[15] , \A_DOUT_TEMPR60[15] , 
        \A_DOUT_TEMPR61[15] , \A_DOUT_TEMPR62[15] , 
        \A_DOUT_TEMPR63[15] , \A_DOUT_TEMPR64[15] , 
        \A_DOUT_TEMPR65[15] , \A_DOUT_TEMPR66[15] , 
        \A_DOUT_TEMPR67[15] , \A_DOUT_TEMPR68[15] , 
        \A_DOUT_TEMPR69[15] , \A_DOUT_TEMPR70[15] , 
        \A_DOUT_TEMPR71[15] , \A_DOUT_TEMPR72[15] , 
        \A_DOUT_TEMPR73[15] , \A_DOUT_TEMPR74[15] , 
        \A_DOUT_TEMPR75[15] , \A_DOUT_TEMPR76[15] , 
        \A_DOUT_TEMPR77[15] , \A_DOUT_TEMPR78[15] , 
        \A_DOUT_TEMPR79[15] , \A_DOUT_TEMPR80[15] , 
        \A_DOUT_TEMPR81[15] , \A_DOUT_TEMPR82[15] , 
        \A_DOUT_TEMPR83[15] , \A_DOUT_TEMPR84[15] , 
        \A_DOUT_TEMPR85[15] , \A_DOUT_TEMPR86[15] , 
        \A_DOUT_TEMPR87[15] , \A_DOUT_TEMPR88[15] , 
        \A_DOUT_TEMPR89[15] , \A_DOUT_TEMPR90[15] , 
        \A_DOUT_TEMPR91[15] , \A_DOUT_TEMPR92[15] , 
        \A_DOUT_TEMPR93[15] , \A_DOUT_TEMPR94[15] , 
        \A_DOUT_TEMPR95[15] , \A_DOUT_TEMPR96[15] , 
        \A_DOUT_TEMPR97[15] , \A_DOUT_TEMPR98[15] , 
        \A_DOUT_TEMPR99[15] , \A_DOUT_TEMPR100[15] , 
        \A_DOUT_TEMPR101[15] , \A_DOUT_TEMPR102[15] , 
        \A_DOUT_TEMPR103[15] , \A_DOUT_TEMPR104[15] , 
        \A_DOUT_TEMPR105[15] , \A_DOUT_TEMPR106[15] , 
        \A_DOUT_TEMPR107[15] , \A_DOUT_TEMPR108[15] , 
        \A_DOUT_TEMPR109[15] , \A_DOUT_TEMPR110[15] , 
        \A_DOUT_TEMPR111[15] , \A_DOUT_TEMPR112[15] , 
        \A_DOUT_TEMPR113[15] , \A_DOUT_TEMPR114[15] , 
        \A_DOUT_TEMPR115[15] , \A_DOUT_TEMPR116[15] , 
        \A_DOUT_TEMPR117[15] , \A_DOUT_TEMPR118[15] , 
        \A_DOUT_TEMPR0[16] , \A_DOUT_TEMPR1[16] , \A_DOUT_TEMPR2[16] , 
        \A_DOUT_TEMPR3[16] , \A_DOUT_TEMPR4[16] , \A_DOUT_TEMPR5[16] , 
        \A_DOUT_TEMPR6[16] , \A_DOUT_TEMPR7[16] , \A_DOUT_TEMPR8[16] , 
        \A_DOUT_TEMPR9[16] , \A_DOUT_TEMPR10[16] , 
        \A_DOUT_TEMPR11[16] , \A_DOUT_TEMPR12[16] , 
        \A_DOUT_TEMPR13[16] , \A_DOUT_TEMPR14[16] , 
        \A_DOUT_TEMPR15[16] , \A_DOUT_TEMPR16[16] , 
        \A_DOUT_TEMPR17[16] , \A_DOUT_TEMPR18[16] , 
        \A_DOUT_TEMPR19[16] , \A_DOUT_TEMPR20[16] , 
        \A_DOUT_TEMPR21[16] , \A_DOUT_TEMPR22[16] , 
        \A_DOUT_TEMPR23[16] , \A_DOUT_TEMPR24[16] , 
        \A_DOUT_TEMPR25[16] , \A_DOUT_TEMPR26[16] , 
        \A_DOUT_TEMPR27[16] , \A_DOUT_TEMPR28[16] , 
        \A_DOUT_TEMPR29[16] , \A_DOUT_TEMPR30[16] , 
        \A_DOUT_TEMPR31[16] , \A_DOUT_TEMPR32[16] , 
        \A_DOUT_TEMPR33[16] , \A_DOUT_TEMPR34[16] , 
        \A_DOUT_TEMPR35[16] , \A_DOUT_TEMPR36[16] , 
        \A_DOUT_TEMPR37[16] , \A_DOUT_TEMPR38[16] , 
        \A_DOUT_TEMPR39[16] , \A_DOUT_TEMPR40[16] , 
        \A_DOUT_TEMPR41[16] , \A_DOUT_TEMPR42[16] , 
        \A_DOUT_TEMPR43[16] , \A_DOUT_TEMPR44[16] , 
        \A_DOUT_TEMPR45[16] , \A_DOUT_TEMPR46[16] , 
        \A_DOUT_TEMPR47[16] , \A_DOUT_TEMPR48[16] , 
        \A_DOUT_TEMPR49[16] , \A_DOUT_TEMPR50[16] , 
        \A_DOUT_TEMPR51[16] , \A_DOUT_TEMPR52[16] , 
        \A_DOUT_TEMPR53[16] , \A_DOUT_TEMPR54[16] , 
        \A_DOUT_TEMPR55[16] , \A_DOUT_TEMPR56[16] , 
        \A_DOUT_TEMPR57[16] , \A_DOUT_TEMPR58[16] , 
        \A_DOUT_TEMPR59[16] , \A_DOUT_TEMPR60[16] , 
        \A_DOUT_TEMPR61[16] , \A_DOUT_TEMPR62[16] , 
        \A_DOUT_TEMPR63[16] , \A_DOUT_TEMPR64[16] , 
        \A_DOUT_TEMPR65[16] , \A_DOUT_TEMPR66[16] , 
        \A_DOUT_TEMPR67[16] , \A_DOUT_TEMPR68[16] , 
        \A_DOUT_TEMPR69[16] , \A_DOUT_TEMPR70[16] , 
        \A_DOUT_TEMPR71[16] , \A_DOUT_TEMPR72[16] , 
        \A_DOUT_TEMPR73[16] , \A_DOUT_TEMPR74[16] , 
        \A_DOUT_TEMPR75[16] , \A_DOUT_TEMPR76[16] , 
        \A_DOUT_TEMPR77[16] , \A_DOUT_TEMPR78[16] , 
        \A_DOUT_TEMPR79[16] , \A_DOUT_TEMPR80[16] , 
        \A_DOUT_TEMPR81[16] , \A_DOUT_TEMPR82[16] , 
        \A_DOUT_TEMPR83[16] , \A_DOUT_TEMPR84[16] , 
        \A_DOUT_TEMPR85[16] , \A_DOUT_TEMPR86[16] , 
        \A_DOUT_TEMPR87[16] , \A_DOUT_TEMPR88[16] , 
        \A_DOUT_TEMPR89[16] , \A_DOUT_TEMPR90[16] , 
        \A_DOUT_TEMPR91[16] , \A_DOUT_TEMPR92[16] , 
        \A_DOUT_TEMPR93[16] , \A_DOUT_TEMPR94[16] , 
        \A_DOUT_TEMPR95[16] , \A_DOUT_TEMPR96[16] , 
        \A_DOUT_TEMPR97[16] , \A_DOUT_TEMPR98[16] , 
        \A_DOUT_TEMPR99[16] , \A_DOUT_TEMPR100[16] , 
        \A_DOUT_TEMPR101[16] , \A_DOUT_TEMPR102[16] , 
        \A_DOUT_TEMPR103[16] , \A_DOUT_TEMPR104[16] , 
        \A_DOUT_TEMPR105[16] , \A_DOUT_TEMPR106[16] , 
        \A_DOUT_TEMPR107[16] , \A_DOUT_TEMPR108[16] , 
        \A_DOUT_TEMPR109[16] , \A_DOUT_TEMPR110[16] , 
        \A_DOUT_TEMPR111[16] , \A_DOUT_TEMPR112[16] , 
        \A_DOUT_TEMPR113[16] , \A_DOUT_TEMPR114[16] , 
        \A_DOUT_TEMPR115[16] , \A_DOUT_TEMPR116[16] , 
        \A_DOUT_TEMPR117[16] , \A_DOUT_TEMPR118[16] , 
        \A_DOUT_TEMPR0[17] , \A_DOUT_TEMPR1[17] , \A_DOUT_TEMPR2[17] , 
        \A_DOUT_TEMPR3[17] , \A_DOUT_TEMPR4[17] , \A_DOUT_TEMPR5[17] , 
        \A_DOUT_TEMPR6[17] , \A_DOUT_TEMPR7[17] , \A_DOUT_TEMPR8[17] , 
        \A_DOUT_TEMPR9[17] , \A_DOUT_TEMPR10[17] , 
        \A_DOUT_TEMPR11[17] , \A_DOUT_TEMPR12[17] , 
        \A_DOUT_TEMPR13[17] , \A_DOUT_TEMPR14[17] , 
        \A_DOUT_TEMPR15[17] , \A_DOUT_TEMPR16[17] , 
        \A_DOUT_TEMPR17[17] , \A_DOUT_TEMPR18[17] , 
        \A_DOUT_TEMPR19[17] , \A_DOUT_TEMPR20[17] , 
        \A_DOUT_TEMPR21[17] , \A_DOUT_TEMPR22[17] , 
        \A_DOUT_TEMPR23[17] , \A_DOUT_TEMPR24[17] , 
        \A_DOUT_TEMPR25[17] , \A_DOUT_TEMPR26[17] , 
        \A_DOUT_TEMPR27[17] , \A_DOUT_TEMPR28[17] , 
        \A_DOUT_TEMPR29[17] , \A_DOUT_TEMPR30[17] , 
        \A_DOUT_TEMPR31[17] , \A_DOUT_TEMPR32[17] , 
        \A_DOUT_TEMPR33[17] , \A_DOUT_TEMPR34[17] , 
        \A_DOUT_TEMPR35[17] , \A_DOUT_TEMPR36[17] , 
        \A_DOUT_TEMPR37[17] , \A_DOUT_TEMPR38[17] , 
        \A_DOUT_TEMPR39[17] , \A_DOUT_TEMPR40[17] , 
        \A_DOUT_TEMPR41[17] , \A_DOUT_TEMPR42[17] , 
        \A_DOUT_TEMPR43[17] , \A_DOUT_TEMPR44[17] , 
        \A_DOUT_TEMPR45[17] , \A_DOUT_TEMPR46[17] , 
        \A_DOUT_TEMPR47[17] , \A_DOUT_TEMPR48[17] , 
        \A_DOUT_TEMPR49[17] , \A_DOUT_TEMPR50[17] , 
        \A_DOUT_TEMPR51[17] , \A_DOUT_TEMPR52[17] , 
        \A_DOUT_TEMPR53[17] , \A_DOUT_TEMPR54[17] , 
        \A_DOUT_TEMPR55[17] , \A_DOUT_TEMPR56[17] , 
        \A_DOUT_TEMPR57[17] , \A_DOUT_TEMPR58[17] , 
        \A_DOUT_TEMPR59[17] , \A_DOUT_TEMPR60[17] , 
        \A_DOUT_TEMPR61[17] , \A_DOUT_TEMPR62[17] , 
        \A_DOUT_TEMPR63[17] , \A_DOUT_TEMPR64[17] , 
        \A_DOUT_TEMPR65[17] , \A_DOUT_TEMPR66[17] , 
        \A_DOUT_TEMPR67[17] , \A_DOUT_TEMPR68[17] , 
        \A_DOUT_TEMPR69[17] , \A_DOUT_TEMPR70[17] , 
        \A_DOUT_TEMPR71[17] , \A_DOUT_TEMPR72[17] , 
        \A_DOUT_TEMPR73[17] , \A_DOUT_TEMPR74[17] , 
        \A_DOUT_TEMPR75[17] , \A_DOUT_TEMPR76[17] , 
        \A_DOUT_TEMPR77[17] , \A_DOUT_TEMPR78[17] , 
        \A_DOUT_TEMPR79[17] , \A_DOUT_TEMPR80[17] , 
        \A_DOUT_TEMPR81[17] , \A_DOUT_TEMPR82[17] , 
        \A_DOUT_TEMPR83[17] , \A_DOUT_TEMPR84[17] , 
        \A_DOUT_TEMPR85[17] , \A_DOUT_TEMPR86[17] , 
        \A_DOUT_TEMPR87[17] , \A_DOUT_TEMPR88[17] , 
        \A_DOUT_TEMPR89[17] , \A_DOUT_TEMPR90[17] , 
        \A_DOUT_TEMPR91[17] , \A_DOUT_TEMPR92[17] , 
        \A_DOUT_TEMPR93[17] , \A_DOUT_TEMPR94[17] , 
        \A_DOUT_TEMPR95[17] , \A_DOUT_TEMPR96[17] , 
        \A_DOUT_TEMPR97[17] , \A_DOUT_TEMPR98[17] , 
        \A_DOUT_TEMPR99[17] , \A_DOUT_TEMPR100[17] , 
        \A_DOUT_TEMPR101[17] , \A_DOUT_TEMPR102[17] , 
        \A_DOUT_TEMPR103[17] , \A_DOUT_TEMPR104[17] , 
        \A_DOUT_TEMPR105[17] , \A_DOUT_TEMPR106[17] , 
        \A_DOUT_TEMPR107[17] , \A_DOUT_TEMPR108[17] , 
        \A_DOUT_TEMPR109[17] , \A_DOUT_TEMPR110[17] , 
        \A_DOUT_TEMPR111[17] , \A_DOUT_TEMPR112[17] , 
        \A_DOUT_TEMPR113[17] , \A_DOUT_TEMPR114[17] , 
        \A_DOUT_TEMPR115[17] , \A_DOUT_TEMPR116[17] , 
        \A_DOUT_TEMPR117[17] , \A_DOUT_TEMPR118[17] , 
        \A_DOUT_TEMPR0[18] , \A_DOUT_TEMPR1[18] , \A_DOUT_TEMPR2[18] , 
        \A_DOUT_TEMPR3[18] , \A_DOUT_TEMPR4[18] , \A_DOUT_TEMPR5[18] , 
        \A_DOUT_TEMPR6[18] , \A_DOUT_TEMPR7[18] , \A_DOUT_TEMPR8[18] , 
        \A_DOUT_TEMPR9[18] , \A_DOUT_TEMPR10[18] , 
        \A_DOUT_TEMPR11[18] , \A_DOUT_TEMPR12[18] , 
        \A_DOUT_TEMPR13[18] , \A_DOUT_TEMPR14[18] , 
        \A_DOUT_TEMPR15[18] , \A_DOUT_TEMPR16[18] , 
        \A_DOUT_TEMPR17[18] , \A_DOUT_TEMPR18[18] , 
        \A_DOUT_TEMPR19[18] , \A_DOUT_TEMPR20[18] , 
        \A_DOUT_TEMPR21[18] , \A_DOUT_TEMPR22[18] , 
        \A_DOUT_TEMPR23[18] , \A_DOUT_TEMPR24[18] , 
        \A_DOUT_TEMPR25[18] , \A_DOUT_TEMPR26[18] , 
        \A_DOUT_TEMPR27[18] , \A_DOUT_TEMPR28[18] , 
        \A_DOUT_TEMPR29[18] , \A_DOUT_TEMPR30[18] , 
        \A_DOUT_TEMPR31[18] , \A_DOUT_TEMPR32[18] , 
        \A_DOUT_TEMPR33[18] , \A_DOUT_TEMPR34[18] , 
        \A_DOUT_TEMPR35[18] , \A_DOUT_TEMPR36[18] , 
        \A_DOUT_TEMPR37[18] , \A_DOUT_TEMPR38[18] , 
        \A_DOUT_TEMPR39[18] , \A_DOUT_TEMPR40[18] , 
        \A_DOUT_TEMPR41[18] , \A_DOUT_TEMPR42[18] , 
        \A_DOUT_TEMPR43[18] , \A_DOUT_TEMPR44[18] , 
        \A_DOUT_TEMPR45[18] , \A_DOUT_TEMPR46[18] , 
        \A_DOUT_TEMPR47[18] , \A_DOUT_TEMPR48[18] , 
        \A_DOUT_TEMPR49[18] , \A_DOUT_TEMPR50[18] , 
        \A_DOUT_TEMPR51[18] , \A_DOUT_TEMPR52[18] , 
        \A_DOUT_TEMPR53[18] , \A_DOUT_TEMPR54[18] , 
        \A_DOUT_TEMPR55[18] , \A_DOUT_TEMPR56[18] , 
        \A_DOUT_TEMPR57[18] , \A_DOUT_TEMPR58[18] , 
        \A_DOUT_TEMPR59[18] , \A_DOUT_TEMPR60[18] , 
        \A_DOUT_TEMPR61[18] , \A_DOUT_TEMPR62[18] , 
        \A_DOUT_TEMPR63[18] , \A_DOUT_TEMPR64[18] , 
        \A_DOUT_TEMPR65[18] , \A_DOUT_TEMPR66[18] , 
        \A_DOUT_TEMPR67[18] , \A_DOUT_TEMPR68[18] , 
        \A_DOUT_TEMPR69[18] , \A_DOUT_TEMPR70[18] , 
        \A_DOUT_TEMPR71[18] , \A_DOUT_TEMPR72[18] , 
        \A_DOUT_TEMPR73[18] , \A_DOUT_TEMPR74[18] , 
        \A_DOUT_TEMPR75[18] , \A_DOUT_TEMPR76[18] , 
        \A_DOUT_TEMPR77[18] , \A_DOUT_TEMPR78[18] , 
        \A_DOUT_TEMPR79[18] , \A_DOUT_TEMPR80[18] , 
        \A_DOUT_TEMPR81[18] , \A_DOUT_TEMPR82[18] , 
        \A_DOUT_TEMPR83[18] , \A_DOUT_TEMPR84[18] , 
        \A_DOUT_TEMPR85[18] , \A_DOUT_TEMPR86[18] , 
        \A_DOUT_TEMPR87[18] , \A_DOUT_TEMPR88[18] , 
        \A_DOUT_TEMPR89[18] , \A_DOUT_TEMPR90[18] , 
        \A_DOUT_TEMPR91[18] , \A_DOUT_TEMPR92[18] , 
        \A_DOUT_TEMPR93[18] , \A_DOUT_TEMPR94[18] , 
        \A_DOUT_TEMPR95[18] , \A_DOUT_TEMPR96[18] , 
        \A_DOUT_TEMPR97[18] , \A_DOUT_TEMPR98[18] , 
        \A_DOUT_TEMPR99[18] , \A_DOUT_TEMPR100[18] , 
        \A_DOUT_TEMPR101[18] , \A_DOUT_TEMPR102[18] , 
        \A_DOUT_TEMPR103[18] , \A_DOUT_TEMPR104[18] , 
        \A_DOUT_TEMPR105[18] , \A_DOUT_TEMPR106[18] , 
        \A_DOUT_TEMPR107[18] , \A_DOUT_TEMPR108[18] , 
        \A_DOUT_TEMPR109[18] , \A_DOUT_TEMPR110[18] , 
        \A_DOUT_TEMPR111[18] , \A_DOUT_TEMPR112[18] , 
        \A_DOUT_TEMPR113[18] , \A_DOUT_TEMPR114[18] , 
        \A_DOUT_TEMPR115[18] , \A_DOUT_TEMPR116[18] , 
        \A_DOUT_TEMPR117[18] , \A_DOUT_TEMPR118[18] , 
        \A_DOUT_TEMPR0[19] , \A_DOUT_TEMPR1[19] , \A_DOUT_TEMPR2[19] , 
        \A_DOUT_TEMPR3[19] , \A_DOUT_TEMPR4[19] , \A_DOUT_TEMPR5[19] , 
        \A_DOUT_TEMPR6[19] , \A_DOUT_TEMPR7[19] , \A_DOUT_TEMPR8[19] , 
        \A_DOUT_TEMPR9[19] , \A_DOUT_TEMPR10[19] , 
        \A_DOUT_TEMPR11[19] , \A_DOUT_TEMPR12[19] , 
        \A_DOUT_TEMPR13[19] , \A_DOUT_TEMPR14[19] , 
        \A_DOUT_TEMPR15[19] , \A_DOUT_TEMPR16[19] , 
        \A_DOUT_TEMPR17[19] , \A_DOUT_TEMPR18[19] , 
        \A_DOUT_TEMPR19[19] , \A_DOUT_TEMPR20[19] , 
        \A_DOUT_TEMPR21[19] , \A_DOUT_TEMPR22[19] , 
        \A_DOUT_TEMPR23[19] , \A_DOUT_TEMPR24[19] , 
        \A_DOUT_TEMPR25[19] , \A_DOUT_TEMPR26[19] , 
        \A_DOUT_TEMPR27[19] , \A_DOUT_TEMPR28[19] , 
        \A_DOUT_TEMPR29[19] , \A_DOUT_TEMPR30[19] , 
        \A_DOUT_TEMPR31[19] , \A_DOUT_TEMPR32[19] , 
        \A_DOUT_TEMPR33[19] , \A_DOUT_TEMPR34[19] , 
        \A_DOUT_TEMPR35[19] , \A_DOUT_TEMPR36[19] , 
        \A_DOUT_TEMPR37[19] , \A_DOUT_TEMPR38[19] , 
        \A_DOUT_TEMPR39[19] , \A_DOUT_TEMPR40[19] , 
        \A_DOUT_TEMPR41[19] , \A_DOUT_TEMPR42[19] , 
        \A_DOUT_TEMPR43[19] , \A_DOUT_TEMPR44[19] , 
        \A_DOUT_TEMPR45[19] , \A_DOUT_TEMPR46[19] , 
        \A_DOUT_TEMPR47[19] , \A_DOUT_TEMPR48[19] , 
        \A_DOUT_TEMPR49[19] , \A_DOUT_TEMPR50[19] , 
        \A_DOUT_TEMPR51[19] , \A_DOUT_TEMPR52[19] , 
        \A_DOUT_TEMPR53[19] , \A_DOUT_TEMPR54[19] , 
        \A_DOUT_TEMPR55[19] , \A_DOUT_TEMPR56[19] , 
        \A_DOUT_TEMPR57[19] , \A_DOUT_TEMPR58[19] , 
        \A_DOUT_TEMPR59[19] , \A_DOUT_TEMPR60[19] , 
        \A_DOUT_TEMPR61[19] , \A_DOUT_TEMPR62[19] , 
        \A_DOUT_TEMPR63[19] , \A_DOUT_TEMPR64[19] , 
        \A_DOUT_TEMPR65[19] , \A_DOUT_TEMPR66[19] , 
        \A_DOUT_TEMPR67[19] , \A_DOUT_TEMPR68[19] , 
        \A_DOUT_TEMPR69[19] , \A_DOUT_TEMPR70[19] , 
        \A_DOUT_TEMPR71[19] , \A_DOUT_TEMPR72[19] , 
        \A_DOUT_TEMPR73[19] , \A_DOUT_TEMPR74[19] , 
        \A_DOUT_TEMPR75[19] , \A_DOUT_TEMPR76[19] , 
        \A_DOUT_TEMPR77[19] , \A_DOUT_TEMPR78[19] , 
        \A_DOUT_TEMPR79[19] , \A_DOUT_TEMPR80[19] , 
        \A_DOUT_TEMPR81[19] , \A_DOUT_TEMPR82[19] , 
        \A_DOUT_TEMPR83[19] , \A_DOUT_TEMPR84[19] , 
        \A_DOUT_TEMPR85[19] , \A_DOUT_TEMPR86[19] , 
        \A_DOUT_TEMPR87[19] , \A_DOUT_TEMPR88[19] , 
        \A_DOUT_TEMPR89[19] , \A_DOUT_TEMPR90[19] , 
        \A_DOUT_TEMPR91[19] , \A_DOUT_TEMPR92[19] , 
        \A_DOUT_TEMPR93[19] , \A_DOUT_TEMPR94[19] , 
        \A_DOUT_TEMPR95[19] , \A_DOUT_TEMPR96[19] , 
        \A_DOUT_TEMPR97[19] , \A_DOUT_TEMPR98[19] , 
        \A_DOUT_TEMPR99[19] , \A_DOUT_TEMPR100[19] , 
        \A_DOUT_TEMPR101[19] , \A_DOUT_TEMPR102[19] , 
        \A_DOUT_TEMPR103[19] , \A_DOUT_TEMPR104[19] , 
        \A_DOUT_TEMPR105[19] , \A_DOUT_TEMPR106[19] , 
        \A_DOUT_TEMPR107[19] , \A_DOUT_TEMPR108[19] , 
        \A_DOUT_TEMPR109[19] , \A_DOUT_TEMPR110[19] , 
        \A_DOUT_TEMPR111[19] , \A_DOUT_TEMPR112[19] , 
        \A_DOUT_TEMPR113[19] , \A_DOUT_TEMPR114[19] , 
        \A_DOUT_TEMPR115[19] , \A_DOUT_TEMPR116[19] , 
        \A_DOUT_TEMPR117[19] , \A_DOUT_TEMPR118[19] , 
        \A_DOUT_TEMPR0[20] , \A_DOUT_TEMPR1[20] , \A_DOUT_TEMPR2[20] , 
        \A_DOUT_TEMPR3[20] , \A_DOUT_TEMPR4[20] , \A_DOUT_TEMPR5[20] , 
        \A_DOUT_TEMPR6[20] , \A_DOUT_TEMPR7[20] , \A_DOUT_TEMPR8[20] , 
        \A_DOUT_TEMPR9[20] , \A_DOUT_TEMPR10[20] , 
        \A_DOUT_TEMPR11[20] , \A_DOUT_TEMPR12[20] , 
        \A_DOUT_TEMPR13[20] , \A_DOUT_TEMPR14[20] , 
        \A_DOUT_TEMPR15[20] , \A_DOUT_TEMPR16[20] , 
        \A_DOUT_TEMPR17[20] , \A_DOUT_TEMPR18[20] , 
        \A_DOUT_TEMPR19[20] , \A_DOUT_TEMPR20[20] , 
        \A_DOUT_TEMPR21[20] , \A_DOUT_TEMPR22[20] , 
        \A_DOUT_TEMPR23[20] , \A_DOUT_TEMPR24[20] , 
        \A_DOUT_TEMPR25[20] , \A_DOUT_TEMPR26[20] , 
        \A_DOUT_TEMPR27[20] , \A_DOUT_TEMPR28[20] , 
        \A_DOUT_TEMPR29[20] , \A_DOUT_TEMPR30[20] , 
        \A_DOUT_TEMPR31[20] , \A_DOUT_TEMPR32[20] , 
        \A_DOUT_TEMPR33[20] , \A_DOUT_TEMPR34[20] , 
        \A_DOUT_TEMPR35[20] , \A_DOUT_TEMPR36[20] , 
        \A_DOUT_TEMPR37[20] , \A_DOUT_TEMPR38[20] , 
        \A_DOUT_TEMPR39[20] , \A_DOUT_TEMPR40[20] , 
        \A_DOUT_TEMPR41[20] , \A_DOUT_TEMPR42[20] , 
        \A_DOUT_TEMPR43[20] , \A_DOUT_TEMPR44[20] , 
        \A_DOUT_TEMPR45[20] , \A_DOUT_TEMPR46[20] , 
        \A_DOUT_TEMPR47[20] , \A_DOUT_TEMPR48[20] , 
        \A_DOUT_TEMPR49[20] , \A_DOUT_TEMPR50[20] , 
        \A_DOUT_TEMPR51[20] , \A_DOUT_TEMPR52[20] , 
        \A_DOUT_TEMPR53[20] , \A_DOUT_TEMPR54[20] , 
        \A_DOUT_TEMPR55[20] , \A_DOUT_TEMPR56[20] , 
        \A_DOUT_TEMPR57[20] , \A_DOUT_TEMPR58[20] , 
        \A_DOUT_TEMPR59[20] , \A_DOUT_TEMPR60[20] , 
        \A_DOUT_TEMPR61[20] , \A_DOUT_TEMPR62[20] , 
        \A_DOUT_TEMPR63[20] , \A_DOUT_TEMPR64[20] , 
        \A_DOUT_TEMPR65[20] , \A_DOUT_TEMPR66[20] , 
        \A_DOUT_TEMPR67[20] , \A_DOUT_TEMPR68[20] , 
        \A_DOUT_TEMPR69[20] , \A_DOUT_TEMPR70[20] , 
        \A_DOUT_TEMPR71[20] , \A_DOUT_TEMPR72[20] , 
        \A_DOUT_TEMPR73[20] , \A_DOUT_TEMPR74[20] , 
        \A_DOUT_TEMPR75[20] , \A_DOUT_TEMPR76[20] , 
        \A_DOUT_TEMPR77[20] , \A_DOUT_TEMPR78[20] , 
        \A_DOUT_TEMPR79[20] , \A_DOUT_TEMPR80[20] , 
        \A_DOUT_TEMPR81[20] , \A_DOUT_TEMPR82[20] , 
        \A_DOUT_TEMPR83[20] , \A_DOUT_TEMPR84[20] , 
        \A_DOUT_TEMPR85[20] , \A_DOUT_TEMPR86[20] , 
        \A_DOUT_TEMPR87[20] , \A_DOUT_TEMPR88[20] , 
        \A_DOUT_TEMPR89[20] , \A_DOUT_TEMPR90[20] , 
        \A_DOUT_TEMPR91[20] , \A_DOUT_TEMPR92[20] , 
        \A_DOUT_TEMPR93[20] , \A_DOUT_TEMPR94[20] , 
        \A_DOUT_TEMPR95[20] , \A_DOUT_TEMPR96[20] , 
        \A_DOUT_TEMPR97[20] , \A_DOUT_TEMPR98[20] , 
        \A_DOUT_TEMPR99[20] , \A_DOUT_TEMPR100[20] , 
        \A_DOUT_TEMPR101[20] , \A_DOUT_TEMPR102[20] , 
        \A_DOUT_TEMPR103[20] , \A_DOUT_TEMPR104[20] , 
        \A_DOUT_TEMPR105[20] , \A_DOUT_TEMPR106[20] , 
        \A_DOUT_TEMPR107[20] , \A_DOUT_TEMPR108[20] , 
        \A_DOUT_TEMPR109[20] , \A_DOUT_TEMPR110[20] , 
        \A_DOUT_TEMPR111[20] , \A_DOUT_TEMPR112[20] , 
        \A_DOUT_TEMPR113[20] , \A_DOUT_TEMPR114[20] , 
        \A_DOUT_TEMPR115[20] , \A_DOUT_TEMPR116[20] , 
        \A_DOUT_TEMPR117[20] , \A_DOUT_TEMPR118[20] , 
        \A_DOUT_TEMPR0[21] , \A_DOUT_TEMPR1[21] , \A_DOUT_TEMPR2[21] , 
        \A_DOUT_TEMPR3[21] , \A_DOUT_TEMPR4[21] , \A_DOUT_TEMPR5[21] , 
        \A_DOUT_TEMPR6[21] , \A_DOUT_TEMPR7[21] , \A_DOUT_TEMPR8[21] , 
        \A_DOUT_TEMPR9[21] , \A_DOUT_TEMPR10[21] , 
        \A_DOUT_TEMPR11[21] , \A_DOUT_TEMPR12[21] , 
        \A_DOUT_TEMPR13[21] , \A_DOUT_TEMPR14[21] , 
        \A_DOUT_TEMPR15[21] , \A_DOUT_TEMPR16[21] , 
        \A_DOUT_TEMPR17[21] , \A_DOUT_TEMPR18[21] , 
        \A_DOUT_TEMPR19[21] , \A_DOUT_TEMPR20[21] , 
        \A_DOUT_TEMPR21[21] , \A_DOUT_TEMPR22[21] , 
        \A_DOUT_TEMPR23[21] , \A_DOUT_TEMPR24[21] , 
        \A_DOUT_TEMPR25[21] , \A_DOUT_TEMPR26[21] , 
        \A_DOUT_TEMPR27[21] , \A_DOUT_TEMPR28[21] , 
        \A_DOUT_TEMPR29[21] , \A_DOUT_TEMPR30[21] , 
        \A_DOUT_TEMPR31[21] , \A_DOUT_TEMPR32[21] , 
        \A_DOUT_TEMPR33[21] , \A_DOUT_TEMPR34[21] , 
        \A_DOUT_TEMPR35[21] , \A_DOUT_TEMPR36[21] , 
        \A_DOUT_TEMPR37[21] , \A_DOUT_TEMPR38[21] , 
        \A_DOUT_TEMPR39[21] , \A_DOUT_TEMPR40[21] , 
        \A_DOUT_TEMPR41[21] , \A_DOUT_TEMPR42[21] , 
        \A_DOUT_TEMPR43[21] , \A_DOUT_TEMPR44[21] , 
        \A_DOUT_TEMPR45[21] , \A_DOUT_TEMPR46[21] , 
        \A_DOUT_TEMPR47[21] , \A_DOUT_TEMPR48[21] , 
        \A_DOUT_TEMPR49[21] , \A_DOUT_TEMPR50[21] , 
        \A_DOUT_TEMPR51[21] , \A_DOUT_TEMPR52[21] , 
        \A_DOUT_TEMPR53[21] , \A_DOUT_TEMPR54[21] , 
        \A_DOUT_TEMPR55[21] , \A_DOUT_TEMPR56[21] , 
        \A_DOUT_TEMPR57[21] , \A_DOUT_TEMPR58[21] , 
        \A_DOUT_TEMPR59[21] , \A_DOUT_TEMPR60[21] , 
        \A_DOUT_TEMPR61[21] , \A_DOUT_TEMPR62[21] , 
        \A_DOUT_TEMPR63[21] , \A_DOUT_TEMPR64[21] , 
        \A_DOUT_TEMPR65[21] , \A_DOUT_TEMPR66[21] , 
        \A_DOUT_TEMPR67[21] , \A_DOUT_TEMPR68[21] , 
        \A_DOUT_TEMPR69[21] , \A_DOUT_TEMPR70[21] , 
        \A_DOUT_TEMPR71[21] , \A_DOUT_TEMPR72[21] , 
        \A_DOUT_TEMPR73[21] , \A_DOUT_TEMPR74[21] , 
        \A_DOUT_TEMPR75[21] , \A_DOUT_TEMPR76[21] , 
        \A_DOUT_TEMPR77[21] , \A_DOUT_TEMPR78[21] , 
        \A_DOUT_TEMPR79[21] , \A_DOUT_TEMPR80[21] , 
        \A_DOUT_TEMPR81[21] , \A_DOUT_TEMPR82[21] , 
        \A_DOUT_TEMPR83[21] , \A_DOUT_TEMPR84[21] , 
        \A_DOUT_TEMPR85[21] , \A_DOUT_TEMPR86[21] , 
        \A_DOUT_TEMPR87[21] , \A_DOUT_TEMPR88[21] , 
        \A_DOUT_TEMPR89[21] , \A_DOUT_TEMPR90[21] , 
        \A_DOUT_TEMPR91[21] , \A_DOUT_TEMPR92[21] , 
        \A_DOUT_TEMPR93[21] , \A_DOUT_TEMPR94[21] , 
        \A_DOUT_TEMPR95[21] , \A_DOUT_TEMPR96[21] , 
        \A_DOUT_TEMPR97[21] , \A_DOUT_TEMPR98[21] , 
        \A_DOUT_TEMPR99[21] , \A_DOUT_TEMPR100[21] , 
        \A_DOUT_TEMPR101[21] , \A_DOUT_TEMPR102[21] , 
        \A_DOUT_TEMPR103[21] , \A_DOUT_TEMPR104[21] , 
        \A_DOUT_TEMPR105[21] , \A_DOUT_TEMPR106[21] , 
        \A_DOUT_TEMPR107[21] , \A_DOUT_TEMPR108[21] , 
        \A_DOUT_TEMPR109[21] , \A_DOUT_TEMPR110[21] , 
        \A_DOUT_TEMPR111[21] , \A_DOUT_TEMPR112[21] , 
        \A_DOUT_TEMPR113[21] , \A_DOUT_TEMPR114[21] , 
        \A_DOUT_TEMPR115[21] , \A_DOUT_TEMPR116[21] , 
        \A_DOUT_TEMPR117[21] , \A_DOUT_TEMPR118[21] , 
        \A_DOUT_TEMPR0[22] , \A_DOUT_TEMPR1[22] , \A_DOUT_TEMPR2[22] , 
        \A_DOUT_TEMPR3[22] , \A_DOUT_TEMPR4[22] , \A_DOUT_TEMPR5[22] , 
        \A_DOUT_TEMPR6[22] , \A_DOUT_TEMPR7[22] , \A_DOUT_TEMPR8[22] , 
        \A_DOUT_TEMPR9[22] , \A_DOUT_TEMPR10[22] , 
        \A_DOUT_TEMPR11[22] , \A_DOUT_TEMPR12[22] , 
        \A_DOUT_TEMPR13[22] , \A_DOUT_TEMPR14[22] , 
        \A_DOUT_TEMPR15[22] , \A_DOUT_TEMPR16[22] , 
        \A_DOUT_TEMPR17[22] , \A_DOUT_TEMPR18[22] , 
        \A_DOUT_TEMPR19[22] , \A_DOUT_TEMPR20[22] , 
        \A_DOUT_TEMPR21[22] , \A_DOUT_TEMPR22[22] , 
        \A_DOUT_TEMPR23[22] , \A_DOUT_TEMPR24[22] , 
        \A_DOUT_TEMPR25[22] , \A_DOUT_TEMPR26[22] , 
        \A_DOUT_TEMPR27[22] , \A_DOUT_TEMPR28[22] , 
        \A_DOUT_TEMPR29[22] , \A_DOUT_TEMPR30[22] , 
        \A_DOUT_TEMPR31[22] , \A_DOUT_TEMPR32[22] , 
        \A_DOUT_TEMPR33[22] , \A_DOUT_TEMPR34[22] , 
        \A_DOUT_TEMPR35[22] , \A_DOUT_TEMPR36[22] , 
        \A_DOUT_TEMPR37[22] , \A_DOUT_TEMPR38[22] , 
        \A_DOUT_TEMPR39[22] , \A_DOUT_TEMPR40[22] , 
        \A_DOUT_TEMPR41[22] , \A_DOUT_TEMPR42[22] , 
        \A_DOUT_TEMPR43[22] , \A_DOUT_TEMPR44[22] , 
        \A_DOUT_TEMPR45[22] , \A_DOUT_TEMPR46[22] , 
        \A_DOUT_TEMPR47[22] , \A_DOUT_TEMPR48[22] , 
        \A_DOUT_TEMPR49[22] , \A_DOUT_TEMPR50[22] , 
        \A_DOUT_TEMPR51[22] , \A_DOUT_TEMPR52[22] , 
        \A_DOUT_TEMPR53[22] , \A_DOUT_TEMPR54[22] , 
        \A_DOUT_TEMPR55[22] , \A_DOUT_TEMPR56[22] , 
        \A_DOUT_TEMPR57[22] , \A_DOUT_TEMPR58[22] , 
        \A_DOUT_TEMPR59[22] , \A_DOUT_TEMPR60[22] , 
        \A_DOUT_TEMPR61[22] , \A_DOUT_TEMPR62[22] , 
        \A_DOUT_TEMPR63[22] , \A_DOUT_TEMPR64[22] , 
        \A_DOUT_TEMPR65[22] , \A_DOUT_TEMPR66[22] , 
        \A_DOUT_TEMPR67[22] , \A_DOUT_TEMPR68[22] , 
        \A_DOUT_TEMPR69[22] , \A_DOUT_TEMPR70[22] , 
        \A_DOUT_TEMPR71[22] , \A_DOUT_TEMPR72[22] , 
        \A_DOUT_TEMPR73[22] , \A_DOUT_TEMPR74[22] , 
        \A_DOUT_TEMPR75[22] , \A_DOUT_TEMPR76[22] , 
        \A_DOUT_TEMPR77[22] , \A_DOUT_TEMPR78[22] , 
        \A_DOUT_TEMPR79[22] , \A_DOUT_TEMPR80[22] , 
        \A_DOUT_TEMPR81[22] , \A_DOUT_TEMPR82[22] , 
        \A_DOUT_TEMPR83[22] , \A_DOUT_TEMPR84[22] , 
        \A_DOUT_TEMPR85[22] , \A_DOUT_TEMPR86[22] , 
        \A_DOUT_TEMPR87[22] , \A_DOUT_TEMPR88[22] , 
        \A_DOUT_TEMPR89[22] , \A_DOUT_TEMPR90[22] , 
        \A_DOUT_TEMPR91[22] , \A_DOUT_TEMPR92[22] , 
        \A_DOUT_TEMPR93[22] , \A_DOUT_TEMPR94[22] , 
        \A_DOUT_TEMPR95[22] , \A_DOUT_TEMPR96[22] , 
        \A_DOUT_TEMPR97[22] , \A_DOUT_TEMPR98[22] , 
        \A_DOUT_TEMPR99[22] , \A_DOUT_TEMPR100[22] , 
        \A_DOUT_TEMPR101[22] , \A_DOUT_TEMPR102[22] , 
        \A_DOUT_TEMPR103[22] , \A_DOUT_TEMPR104[22] , 
        \A_DOUT_TEMPR105[22] , \A_DOUT_TEMPR106[22] , 
        \A_DOUT_TEMPR107[22] , \A_DOUT_TEMPR108[22] , 
        \A_DOUT_TEMPR109[22] , \A_DOUT_TEMPR110[22] , 
        \A_DOUT_TEMPR111[22] , \A_DOUT_TEMPR112[22] , 
        \A_DOUT_TEMPR113[22] , \A_DOUT_TEMPR114[22] , 
        \A_DOUT_TEMPR115[22] , \A_DOUT_TEMPR116[22] , 
        \A_DOUT_TEMPR117[22] , \A_DOUT_TEMPR118[22] , 
        \A_DOUT_TEMPR0[23] , \A_DOUT_TEMPR1[23] , \A_DOUT_TEMPR2[23] , 
        \A_DOUT_TEMPR3[23] , \A_DOUT_TEMPR4[23] , \A_DOUT_TEMPR5[23] , 
        \A_DOUT_TEMPR6[23] , \A_DOUT_TEMPR7[23] , \A_DOUT_TEMPR8[23] , 
        \A_DOUT_TEMPR9[23] , \A_DOUT_TEMPR10[23] , 
        \A_DOUT_TEMPR11[23] , \A_DOUT_TEMPR12[23] , 
        \A_DOUT_TEMPR13[23] , \A_DOUT_TEMPR14[23] , 
        \A_DOUT_TEMPR15[23] , \A_DOUT_TEMPR16[23] , 
        \A_DOUT_TEMPR17[23] , \A_DOUT_TEMPR18[23] , 
        \A_DOUT_TEMPR19[23] , \A_DOUT_TEMPR20[23] , 
        \A_DOUT_TEMPR21[23] , \A_DOUT_TEMPR22[23] , 
        \A_DOUT_TEMPR23[23] , \A_DOUT_TEMPR24[23] , 
        \A_DOUT_TEMPR25[23] , \A_DOUT_TEMPR26[23] , 
        \A_DOUT_TEMPR27[23] , \A_DOUT_TEMPR28[23] , 
        \A_DOUT_TEMPR29[23] , \A_DOUT_TEMPR30[23] , 
        \A_DOUT_TEMPR31[23] , \A_DOUT_TEMPR32[23] , 
        \A_DOUT_TEMPR33[23] , \A_DOUT_TEMPR34[23] , 
        \A_DOUT_TEMPR35[23] , \A_DOUT_TEMPR36[23] , 
        \A_DOUT_TEMPR37[23] , \A_DOUT_TEMPR38[23] , 
        \A_DOUT_TEMPR39[23] , \A_DOUT_TEMPR40[23] , 
        \A_DOUT_TEMPR41[23] , \A_DOUT_TEMPR42[23] , 
        \A_DOUT_TEMPR43[23] , \A_DOUT_TEMPR44[23] , 
        \A_DOUT_TEMPR45[23] , \A_DOUT_TEMPR46[23] , 
        \A_DOUT_TEMPR47[23] , \A_DOUT_TEMPR48[23] , 
        \A_DOUT_TEMPR49[23] , \A_DOUT_TEMPR50[23] , 
        \A_DOUT_TEMPR51[23] , \A_DOUT_TEMPR52[23] , 
        \A_DOUT_TEMPR53[23] , \A_DOUT_TEMPR54[23] , 
        \A_DOUT_TEMPR55[23] , \A_DOUT_TEMPR56[23] , 
        \A_DOUT_TEMPR57[23] , \A_DOUT_TEMPR58[23] , 
        \A_DOUT_TEMPR59[23] , \A_DOUT_TEMPR60[23] , 
        \A_DOUT_TEMPR61[23] , \A_DOUT_TEMPR62[23] , 
        \A_DOUT_TEMPR63[23] , \A_DOUT_TEMPR64[23] , 
        \A_DOUT_TEMPR65[23] , \A_DOUT_TEMPR66[23] , 
        \A_DOUT_TEMPR67[23] , \A_DOUT_TEMPR68[23] , 
        \A_DOUT_TEMPR69[23] , \A_DOUT_TEMPR70[23] , 
        \A_DOUT_TEMPR71[23] , \A_DOUT_TEMPR72[23] , 
        \A_DOUT_TEMPR73[23] , \A_DOUT_TEMPR74[23] , 
        \A_DOUT_TEMPR75[23] , \A_DOUT_TEMPR76[23] , 
        \A_DOUT_TEMPR77[23] , \A_DOUT_TEMPR78[23] , 
        \A_DOUT_TEMPR79[23] , \A_DOUT_TEMPR80[23] , 
        \A_DOUT_TEMPR81[23] , \A_DOUT_TEMPR82[23] , 
        \A_DOUT_TEMPR83[23] , \A_DOUT_TEMPR84[23] , 
        \A_DOUT_TEMPR85[23] , \A_DOUT_TEMPR86[23] , 
        \A_DOUT_TEMPR87[23] , \A_DOUT_TEMPR88[23] , 
        \A_DOUT_TEMPR89[23] , \A_DOUT_TEMPR90[23] , 
        \A_DOUT_TEMPR91[23] , \A_DOUT_TEMPR92[23] , 
        \A_DOUT_TEMPR93[23] , \A_DOUT_TEMPR94[23] , 
        \A_DOUT_TEMPR95[23] , \A_DOUT_TEMPR96[23] , 
        \A_DOUT_TEMPR97[23] , \A_DOUT_TEMPR98[23] , 
        \A_DOUT_TEMPR99[23] , \A_DOUT_TEMPR100[23] , 
        \A_DOUT_TEMPR101[23] , \A_DOUT_TEMPR102[23] , 
        \A_DOUT_TEMPR103[23] , \A_DOUT_TEMPR104[23] , 
        \A_DOUT_TEMPR105[23] , \A_DOUT_TEMPR106[23] , 
        \A_DOUT_TEMPR107[23] , \A_DOUT_TEMPR108[23] , 
        \A_DOUT_TEMPR109[23] , \A_DOUT_TEMPR110[23] , 
        \A_DOUT_TEMPR111[23] , \A_DOUT_TEMPR112[23] , 
        \A_DOUT_TEMPR113[23] , \A_DOUT_TEMPR114[23] , 
        \A_DOUT_TEMPR115[23] , \A_DOUT_TEMPR116[23] , 
        \A_DOUT_TEMPR117[23] , \A_DOUT_TEMPR118[23] , 
        \A_DOUT_TEMPR0[24] , \A_DOUT_TEMPR1[24] , \A_DOUT_TEMPR2[24] , 
        \A_DOUT_TEMPR3[24] , \A_DOUT_TEMPR4[24] , \A_DOUT_TEMPR5[24] , 
        \A_DOUT_TEMPR6[24] , \A_DOUT_TEMPR7[24] , \A_DOUT_TEMPR8[24] , 
        \A_DOUT_TEMPR9[24] , \A_DOUT_TEMPR10[24] , 
        \A_DOUT_TEMPR11[24] , \A_DOUT_TEMPR12[24] , 
        \A_DOUT_TEMPR13[24] , \A_DOUT_TEMPR14[24] , 
        \A_DOUT_TEMPR15[24] , \A_DOUT_TEMPR16[24] , 
        \A_DOUT_TEMPR17[24] , \A_DOUT_TEMPR18[24] , 
        \A_DOUT_TEMPR19[24] , \A_DOUT_TEMPR20[24] , 
        \A_DOUT_TEMPR21[24] , \A_DOUT_TEMPR22[24] , 
        \A_DOUT_TEMPR23[24] , \A_DOUT_TEMPR24[24] , 
        \A_DOUT_TEMPR25[24] , \A_DOUT_TEMPR26[24] , 
        \A_DOUT_TEMPR27[24] , \A_DOUT_TEMPR28[24] , 
        \A_DOUT_TEMPR29[24] , \A_DOUT_TEMPR30[24] , 
        \A_DOUT_TEMPR31[24] , \A_DOUT_TEMPR32[24] , 
        \A_DOUT_TEMPR33[24] , \A_DOUT_TEMPR34[24] , 
        \A_DOUT_TEMPR35[24] , \A_DOUT_TEMPR36[24] , 
        \A_DOUT_TEMPR37[24] , \A_DOUT_TEMPR38[24] , 
        \A_DOUT_TEMPR39[24] , \A_DOUT_TEMPR40[24] , 
        \A_DOUT_TEMPR41[24] , \A_DOUT_TEMPR42[24] , 
        \A_DOUT_TEMPR43[24] , \A_DOUT_TEMPR44[24] , 
        \A_DOUT_TEMPR45[24] , \A_DOUT_TEMPR46[24] , 
        \A_DOUT_TEMPR47[24] , \A_DOUT_TEMPR48[24] , 
        \A_DOUT_TEMPR49[24] , \A_DOUT_TEMPR50[24] , 
        \A_DOUT_TEMPR51[24] , \A_DOUT_TEMPR52[24] , 
        \A_DOUT_TEMPR53[24] , \A_DOUT_TEMPR54[24] , 
        \A_DOUT_TEMPR55[24] , \A_DOUT_TEMPR56[24] , 
        \A_DOUT_TEMPR57[24] , \A_DOUT_TEMPR58[24] , 
        \A_DOUT_TEMPR59[24] , \A_DOUT_TEMPR60[24] , 
        \A_DOUT_TEMPR61[24] , \A_DOUT_TEMPR62[24] , 
        \A_DOUT_TEMPR63[24] , \A_DOUT_TEMPR64[24] , 
        \A_DOUT_TEMPR65[24] , \A_DOUT_TEMPR66[24] , 
        \A_DOUT_TEMPR67[24] , \A_DOUT_TEMPR68[24] , 
        \A_DOUT_TEMPR69[24] , \A_DOUT_TEMPR70[24] , 
        \A_DOUT_TEMPR71[24] , \A_DOUT_TEMPR72[24] , 
        \A_DOUT_TEMPR73[24] , \A_DOUT_TEMPR74[24] , 
        \A_DOUT_TEMPR75[24] , \A_DOUT_TEMPR76[24] , 
        \A_DOUT_TEMPR77[24] , \A_DOUT_TEMPR78[24] , 
        \A_DOUT_TEMPR79[24] , \A_DOUT_TEMPR80[24] , 
        \A_DOUT_TEMPR81[24] , \A_DOUT_TEMPR82[24] , 
        \A_DOUT_TEMPR83[24] , \A_DOUT_TEMPR84[24] , 
        \A_DOUT_TEMPR85[24] , \A_DOUT_TEMPR86[24] , 
        \A_DOUT_TEMPR87[24] , \A_DOUT_TEMPR88[24] , 
        \A_DOUT_TEMPR89[24] , \A_DOUT_TEMPR90[24] , 
        \A_DOUT_TEMPR91[24] , \A_DOUT_TEMPR92[24] , 
        \A_DOUT_TEMPR93[24] , \A_DOUT_TEMPR94[24] , 
        \A_DOUT_TEMPR95[24] , \A_DOUT_TEMPR96[24] , 
        \A_DOUT_TEMPR97[24] , \A_DOUT_TEMPR98[24] , 
        \A_DOUT_TEMPR99[24] , \A_DOUT_TEMPR100[24] , 
        \A_DOUT_TEMPR101[24] , \A_DOUT_TEMPR102[24] , 
        \A_DOUT_TEMPR103[24] , \A_DOUT_TEMPR104[24] , 
        \A_DOUT_TEMPR105[24] , \A_DOUT_TEMPR106[24] , 
        \A_DOUT_TEMPR107[24] , \A_DOUT_TEMPR108[24] , 
        \A_DOUT_TEMPR109[24] , \A_DOUT_TEMPR110[24] , 
        \A_DOUT_TEMPR111[24] , \A_DOUT_TEMPR112[24] , 
        \A_DOUT_TEMPR113[24] , \A_DOUT_TEMPR114[24] , 
        \A_DOUT_TEMPR115[24] , \A_DOUT_TEMPR116[24] , 
        \A_DOUT_TEMPR117[24] , \A_DOUT_TEMPR118[24] , 
        \A_DOUT_TEMPR0[25] , \A_DOUT_TEMPR1[25] , \A_DOUT_TEMPR2[25] , 
        \A_DOUT_TEMPR3[25] , \A_DOUT_TEMPR4[25] , \A_DOUT_TEMPR5[25] , 
        \A_DOUT_TEMPR6[25] , \A_DOUT_TEMPR7[25] , \A_DOUT_TEMPR8[25] , 
        \A_DOUT_TEMPR9[25] , \A_DOUT_TEMPR10[25] , 
        \A_DOUT_TEMPR11[25] , \A_DOUT_TEMPR12[25] , 
        \A_DOUT_TEMPR13[25] , \A_DOUT_TEMPR14[25] , 
        \A_DOUT_TEMPR15[25] , \A_DOUT_TEMPR16[25] , 
        \A_DOUT_TEMPR17[25] , \A_DOUT_TEMPR18[25] , 
        \A_DOUT_TEMPR19[25] , \A_DOUT_TEMPR20[25] , 
        \A_DOUT_TEMPR21[25] , \A_DOUT_TEMPR22[25] , 
        \A_DOUT_TEMPR23[25] , \A_DOUT_TEMPR24[25] , 
        \A_DOUT_TEMPR25[25] , \A_DOUT_TEMPR26[25] , 
        \A_DOUT_TEMPR27[25] , \A_DOUT_TEMPR28[25] , 
        \A_DOUT_TEMPR29[25] , \A_DOUT_TEMPR30[25] , 
        \A_DOUT_TEMPR31[25] , \A_DOUT_TEMPR32[25] , 
        \A_DOUT_TEMPR33[25] , \A_DOUT_TEMPR34[25] , 
        \A_DOUT_TEMPR35[25] , \A_DOUT_TEMPR36[25] , 
        \A_DOUT_TEMPR37[25] , \A_DOUT_TEMPR38[25] , 
        \A_DOUT_TEMPR39[25] , \A_DOUT_TEMPR40[25] , 
        \A_DOUT_TEMPR41[25] , \A_DOUT_TEMPR42[25] , 
        \A_DOUT_TEMPR43[25] , \A_DOUT_TEMPR44[25] , 
        \A_DOUT_TEMPR45[25] , \A_DOUT_TEMPR46[25] , 
        \A_DOUT_TEMPR47[25] , \A_DOUT_TEMPR48[25] , 
        \A_DOUT_TEMPR49[25] , \A_DOUT_TEMPR50[25] , 
        \A_DOUT_TEMPR51[25] , \A_DOUT_TEMPR52[25] , 
        \A_DOUT_TEMPR53[25] , \A_DOUT_TEMPR54[25] , 
        \A_DOUT_TEMPR55[25] , \A_DOUT_TEMPR56[25] , 
        \A_DOUT_TEMPR57[25] , \A_DOUT_TEMPR58[25] , 
        \A_DOUT_TEMPR59[25] , \A_DOUT_TEMPR60[25] , 
        \A_DOUT_TEMPR61[25] , \A_DOUT_TEMPR62[25] , 
        \A_DOUT_TEMPR63[25] , \A_DOUT_TEMPR64[25] , 
        \A_DOUT_TEMPR65[25] , \A_DOUT_TEMPR66[25] , 
        \A_DOUT_TEMPR67[25] , \A_DOUT_TEMPR68[25] , 
        \A_DOUT_TEMPR69[25] , \A_DOUT_TEMPR70[25] , 
        \A_DOUT_TEMPR71[25] , \A_DOUT_TEMPR72[25] , 
        \A_DOUT_TEMPR73[25] , \A_DOUT_TEMPR74[25] , 
        \A_DOUT_TEMPR75[25] , \A_DOUT_TEMPR76[25] , 
        \A_DOUT_TEMPR77[25] , \A_DOUT_TEMPR78[25] , 
        \A_DOUT_TEMPR79[25] , \A_DOUT_TEMPR80[25] , 
        \A_DOUT_TEMPR81[25] , \A_DOUT_TEMPR82[25] , 
        \A_DOUT_TEMPR83[25] , \A_DOUT_TEMPR84[25] , 
        \A_DOUT_TEMPR85[25] , \A_DOUT_TEMPR86[25] , 
        \A_DOUT_TEMPR87[25] , \A_DOUT_TEMPR88[25] , 
        \A_DOUT_TEMPR89[25] , \A_DOUT_TEMPR90[25] , 
        \A_DOUT_TEMPR91[25] , \A_DOUT_TEMPR92[25] , 
        \A_DOUT_TEMPR93[25] , \A_DOUT_TEMPR94[25] , 
        \A_DOUT_TEMPR95[25] , \A_DOUT_TEMPR96[25] , 
        \A_DOUT_TEMPR97[25] , \A_DOUT_TEMPR98[25] , 
        \A_DOUT_TEMPR99[25] , \A_DOUT_TEMPR100[25] , 
        \A_DOUT_TEMPR101[25] , \A_DOUT_TEMPR102[25] , 
        \A_DOUT_TEMPR103[25] , \A_DOUT_TEMPR104[25] , 
        \A_DOUT_TEMPR105[25] , \A_DOUT_TEMPR106[25] , 
        \A_DOUT_TEMPR107[25] , \A_DOUT_TEMPR108[25] , 
        \A_DOUT_TEMPR109[25] , \A_DOUT_TEMPR110[25] , 
        \A_DOUT_TEMPR111[25] , \A_DOUT_TEMPR112[25] , 
        \A_DOUT_TEMPR113[25] , \A_DOUT_TEMPR114[25] , 
        \A_DOUT_TEMPR115[25] , \A_DOUT_TEMPR116[25] , 
        \A_DOUT_TEMPR117[25] , \A_DOUT_TEMPR118[25] , 
        \A_DOUT_TEMPR0[26] , \A_DOUT_TEMPR1[26] , \A_DOUT_TEMPR2[26] , 
        \A_DOUT_TEMPR3[26] , \A_DOUT_TEMPR4[26] , \A_DOUT_TEMPR5[26] , 
        \A_DOUT_TEMPR6[26] , \A_DOUT_TEMPR7[26] , \A_DOUT_TEMPR8[26] , 
        \A_DOUT_TEMPR9[26] , \A_DOUT_TEMPR10[26] , 
        \A_DOUT_TEMPR11[26] , \A_DOUT_TEMPR12[26] , 
        \A_DOUT_TEMPR13[26] , \A_DOUT_TEMPR14[26] , 
        \A_DOUT_TEMPR15[26] , \A_DOUT_TEMPR16[26] , 
        \A_DOUT_TEMPR17[26] , \A_DOUT_TEMPR18[26] , 
        \A_DOUT_TEMPR19[26] , \A_DOUT_TEMPR20[26] , 
        \A_DOUT_TEMPR21[26] , \A_DOUT_TEMPR22[26] , 
        \A_DOUT_TEMPR23[26] , \A_DOUT_TEMPR24[26] , 
        \A_DOUT_TEMPR25[26] , \A_DOUT_TEMPR26[26] , 
        \A_DOUT_TEMPR27[26] , \A_DOUT_TEMPR28[26] , 
        \A_DOUT_TEMPR29[26] , \A_DOUT_TEMPR30[26] , 
        \A_DOUT_TEMPR31[26] , \A_DOUT_TEMPR32[26] , 
        \A_DOUT_TEMPR33[26] , \A_DOUT_TEMPR34[26] , 
        \A_DOUT_TEMPR35[26] , \A_DOUT_TEMPR36[26] , 
        \A_DOUT_TEMPR37[26] , \A_DOUT_TEMPR38[26] , 
        \A_DOUT_TEMPR39[26] , \A_DOUT_TEMPR40[26] , 
        \A_DOUT_TEMPR41[26] , \A_DOUT_TEMPR42[26] , 
        \A_DOUT_TEMPR43[26] , \A_DOUT_TEMPR44[26] , 
        \A_DOUT_TEMPR45[26] , \A_DOUT_TEMPR46[26] , 
        \A_DOUT_TEMPR47[26] , \A_DOUT_TEMPR48[26] , 
        \A_DOUT_TEMPR49[26] , \A_DOUT_TEMPR50[26] , 
        \A_DOUT_TEMPR51[26] , \A_DOUT_TEMPR52[26] , 
        \A_DOUT_TEMPR53[26] , \A_DOUT_TEMPR54[26] , 
        \A_DOUT_TEMPR55[26] , \A_DOUT_TEMPR56[26] , 
        \A_DOUT_TEMPR57[26] , \A_DOUT_TEMPR58[26] , 
        \A_DOUT_TEMPR59[26] , \A_DOUT_TEMPR60[26] , 
        \A_DOUT_TEMPR61[26] , \A_DOUT_TEMPR62[26] , 
        \A_DOUT_TEMPR63[26] , \A_DOUT_TEMPR64[26] , 
        \A_DOUT_TEMPR65[26] , \A_DOUT_TEMPR66[26] , 
        \A_DOUT_TEMPR67[26] , \A_DOUT_TEMPR68[26] , 
        \A_DOUT_TEMPR69[26] , \A_DOUT_TEMPR70[26] , 
        \A_DOUT_TEMPR71[26] , \A_DOUT_TEMPR72[26] , 
        \A_DOUT_TEMPR73[26] , \A_DOUT_TEMPR74[26] , 
        \A_DOUT_TEMPR75[26] , \A_DOUT_TEMPR76[26] , 
        \A_DOUT_TEMPR77[26] , \A_DOUT_TEMPR78[26] , 
        \A_DOUT_TEMPR79[26] , \A_DOUT_TEMPR80[26] , 
        \A_DOUT_TEMPR81[26] , \A_DOUT_TEMPR82[26] , 
        \A_DOUT_TEMPR83[26] , \A_DOUT_TEMPR84[26] , 
        \A_DOUT_TEMPR85[26] , \A_DOUT_TEMPR86[26] , 
        \A_DOUT_TEMPR87[26] , \A_DOUT_TEMPR88[26] , 
        \A_DOUT_TEMPR89[26] , \A_DOUT_TEMPR90[26] , 
        \A_DOUT_TEMPR91[26] , \A_DOUT_TEMPR92[26] , 
        \A_DOUT_TEMPR93[26] , \A_DOUT_TEMPR94[26] , 
        \A_DOUT_TEMPR95[26] , \A_DOUT_TEMPR96[26] , 
        \A_DOUT_TEMPR97[26] , \A_DOUT_TEMPR98[26] , 
        \A_DOUT_TEMPR99[26] , \A_DOUT_TEMPR100[26] , 
        \A_DOUT_TEMPR101[26] , \A_DOUT_TEMPR102[26] , 
        \A_DOUT_TEMPR103[26] , \A_DOUT_TEMPR104[26] , 
        \A_DOUT_TEMPR105[26] , \A_DOUT_TEMPR106[26] , 
        \A_DOUT_TEMPR107[26] , \A_DOUT_TEMPR108[26] , 
        \A_DOUT_TEMPR109[26] , \A_DOUT_TEMPR110[26] , 
        \A_DOUT_TEMPR111[26] , \A_DOUT_TEMPR112[26] , 
        \A_DOUT_TEMPR113[26] , \A_DOUT_TEMPR114[26] , 
        \A_DOUT_TEMPR115[26] , \A_DOUT_TEMPR116[26] , 
        \A_DOUT_TEMPR117[26] , \A_DOUT_TEMPR118[26] , 
        \A_DOUT_TEMPR0[27] , \A_DOUT_TEMPR1[27] , \A_DOUT_TEMPR2[27] , 
        \A_DOUT_TEMPR3[27] , \A_DOUT_TEMPR4[27] , \A_DOUT_TEMPR5[27] , 
        \A_DOUT_TEMPR6[27] , \A_DOUT_TEMPR7[27] , \A_DOUT_TEMPR8[27] , 
        \A_DOUT_TEMPR9[27] , \A_DOUT_TEMPR10[27] , 
        \A_DOUT_TEMPR11[27] , \A_DOUT_TEMPR12[27] , 
        \A_DOUT_TEMPR13[27] , \A_DOUT_TEMPR14[27] , 
        \A_DOUT_TEMPR15[27] , \A_DOUT_TEMPR16[27] , 
        \A_DOUT_TEMPR17[27] , \A_DOUT_TEMPR18[27] , 
        \A_DOUT_TEMPR19[27] , \A_DOUT_TEMPR20[27] , 
        \A_DOUT_TEMPR21[27] , \A_DOUT_TEMPR22[27] , 
        \A_DOUT_TEMPR23[27] , \A_DOUT_TEMPR24[27] , 
        \A_DOUT_TEMPR25[27] , \A_DOUT_TEMPR26[27] , 
        \A_DOUT_TEMPR27[27] , \A_DOUT_TEMPR28[27] , 
        \A_DOUT_TEMPR29[27] , \A_DOUT_TEMPR30[27] , 
        \A_DOUT_TEMPR31[27] , \A_DOUT_TEMPR32[27] , 
        \A_DOUT_TEMPR33[27] , \A_DOUT_TEMPR34[27] , 
        \A_DOUT_TEMPR35[27] , \A_DOUT_TEMPR36[27] , 
        \A_DOUT_TEMPR37[27] , \A_DOUT_TEMPR38[27] , 
        \A_DOUT_TEMPR39[27] , \A_DOUT_TEMPR40[27] , 
        \A_DOUT_TEMPR41[27] , \A_DOUT_TEMPR42[27] , 
        \A_DOUT_TEMPR43[27] , \A_DOUT_TEMPR44[27] , 
        \A_DOUT_TEMPR45[27] , \A_DOUT_TEMPR46[27] , 
        \A_DOUT_TEMPR47[27] , \A_DOUT_TEMPR48[27] , 
        \A_DOUT_TEMPR49[27] , \A_DOUT_TEMPR50[27] , 
        \A_DOUT_TEMPR51[27] , \A_DOUT_TEMPR52[27] , 
        \A_DOUT_TEMPR53[27] , \A_DOUT_TEMPR54[27] , 
        \A_DOUT_TEMPR55[27] , \A_DOUT_TEMPR56[27] , 
        \A_DOUT_TEMPR57[27] , \A_DOUT_TEMPR58[27] , 
        \A_DOUT_TEMPR59[27] , \A_DOUT_TEMPR60[27] , 
        \A_DOUT_TEMPR61[27] , \A_DOUT_TEMPR62[27] , 
        \A_DOUT_TEMPR63[27] , \A_DOUT_TEMPR64[27] , 
        \A_DOUT_TEMPR65[27] , \A_DOUT_TEMPR66[27] , 
        \A_DOUT_TEMPR67[27] , \A_DOUT_TEMPR68[27] , 
        \A_DOUT_TEMPR69[27] , \A_DOUT_TEMPR70[27] , 
        \A_DOUT_TEMPR71[27] , \A_DOUT_TEMPR72[27] , 
        \A_DOUT_TEMPR73[27] , \A_DOUT_TEMPR74[27] , 
        \A_DOUT_TEMPR75[27] , \A_DOUT_TEMPR76[27] , 
        \A_DOUT_TEMPR77[27] , \A_DOUT_TEMPR78[27] , 
        \A_DOUT_TEMPR79[27] , \A_DOUT_TEMPR80[27] , 
        \A_DOUT_TEMPR81[27] , \A_DOUT_TEMPR82[27] , 
        \A_DOUT_TEMPR83[27] , \A_DOUT_TEMPR84[27] , 
        \A_DOUT_TEMPR85[27] , \A_DOUT_TEMPR86[27] , 
        \A_DOUT_TEMPR87[27] , \A_DOUT_TEMPR88[27] , 
        \A_DOUT_TEMPR89[27] , \A_DOUT_TEMPR90[27] , 
        \A_DOUT_TEMPR91[27] , \A_DOUT_TEMPR92[27] , 
        \A_DOUT_TEMPR93[27] , \A_DOUT_TEMPR94[27] , 
        \A_DOUT_TEMPR95[27] , \A_DOUT_TEMPR96[27] , 
        \A_DOUT_TEMPR97[27] , \A_DOUT_TEMPR98[27] , 
        \A_DOUT_TEMPR99[27] , \A_DOUT_TEMPR100[27] , 
        \A_DOUT_TEMPR101[27] , \A_DOUT_TEMPR102[27] , 
        \A_DOUT_TEMPR103[27] , \A_DOUT_TEMPR104[27] , 
        \A_DOUT_TEMPR105[27] , \A_DOUT_TEMPR106[27] , 
        \A_DOUT_TEMPR107[27] , \A_DOUT_TEMPR108[27] , 
        \A_DOUT_TEMPR109[27] , \A_DOUT_TEMPR110[27] , 
        \A_DOUT_TEMPR111[27] , \A_DOUT_TEMPR112[27] , 
        \A_DOUT_TEMPR113[27] , \A_DOUT_TEMPR114[27] , 
        \A_DOUT_TEMPR115[27] , \A_DOUT_TEMPR116[27] , 
        \A_DOUT_TEMPR117[27] , \A_DOUT_TEMPR118[27] , 
        \A_DOUT_TEMPR0[28] , \A_DOUT_TEMPR1[28] , \A_DOUT_TEMPR2[28] , 
        \A_DOUT_TEMPR3[28] , \A_DOUT_TEMPR4[28] , \A_DOUT_TEMPR5[28] , 
        \A_DOUT_TEMPR6[28] , \A_DOUT_TEMPR7[28] , \A_DOUT_TEMPR8[28] , 
        \A_DOUT_TEMPR9[28] , \A_DOUT_TEMPR10[28] , 
        \A_DOUT_TEMPR11[28] , \A_DOUT_TEMPR12[28] , 
        \A_DOUT_TEMPR13[28] , \A_DOUT_TEMPR14[28] , 
        \A_DOUT_TEMPR15[28] , \A_DOUT_TEMPR16[28] , 
        \A_DOUT_TEMPR17[28] , \A_DOUT_TEMPR18[28] , 
        \A_DOUT_TEMPR19[28] , \A_DOUT_TEMPR20[28] , 
        \A_DOUT_TEMPR21[28] , \A_DOUT_TEMPR22[28] , 
        \A_DOUT_TEMPR23[28] , \A_DOUT_TEMPR24[28] , 
        \A_DOUT_TEMPR25[28] , \A_DOUT_TEMPR26[28] , 
        \A_DOUT_TEMPR27[28] , \A_DOUT_TEMPR28[28] , 
        \A_DOUT_TEMPR29[28] , \A_DOUT_TEMPR30[28] , 
        \A_DOUT_TEMPR31[28] , \A_DOUT_TEMPR32[28] , 
        \A_DOUT_TEMPR33[28] , \A_DOUT_TEMPR34[28] , 
        \A_DOUT_TEMPR35[28] , \A_DOUT_TEMPR36[28] , 
        \A_DOUT_TEMPR37[28] , \A_DOUT_TEMPR38[28] , 
        \A_DOUT_TEMPR39[28] , \A_DOUT_TEMPR40[28] , 
        \A_DOUT_TEMPR41[28] , \A_DOUT_TEMPR42[28] , 
        \A_DOUT_TEMPR43[28] , \A_DOUT_TEMPR44[28] , 
        \A_DOUT_TEMPR45[28] , \A_DOUT_TEMPR46[28] , 
        \A_DOUT_TEMPR47[28] , \A_DOUT_TEMPR48[28] , 
        \A_DOUT_TEMPR49[28] , \A_DOUT_TEMPR50[28] , 
        \A_DOUT_TEMPR51[28] , \A_DOUT_TEMPR52[28] , 
        \A_DOUT_TEMPR53[28] , \A_DOUT_TEMPR54[28] , 
        \A_DOUT_TEMPR55[28] , \A_DOUT_TEMPR56[28] , 
        \A_DOUT_TEMPR57[28] , \A_DOUT_TEMPR58[28] , 
        \A_DOUT_TEMPR59[28] , \A_DOUT_TEMPR60[28] , 
        \A_DOUT_TEMPR61[28] , \A_DOUT_TEMPR62[28] , 
        \A_DOUT_TEMPR63[28] , \A_DOUT_TEMPR64[28] , 
        \A_DOUT_TEMPR65[28] , \A_DOUT_TEMPR66[28] , 
        \A_DOUT_TEMPR67[28] , \A_DOUT_TEMPR68[28] , 
        \A_DOUT_TEMPR69[28] , \A_DOUT_TEMPR70[28] , 
        \A_DOUT_TEMPR71[28] , \A_DOUT_TEMPR72[28] , 
        \A_DOUT_TEMPR73[28] , \A_DOUT_TEMPR74[28] , 
        \A_DOUT_TEMPR75[28] , \A_DOUT_TEMPR76[28] , 
        \A_DOUT_TEMPR77[28] , \A_DOUT_TEMPR78[28] , 
        \A_DOUT_TEMPR79[28] , \A_DOUT_TEMPR80[28] , 
        \A_DOUT_TEMPR81[28] , \A_DOUT_TEMPR82[28] , 
        \A_DOUT_TEMPR83[28] , \A_DOUT_TEMPR84[28] , 
        \A_DOUT_TEMPR85[28] , \A_DOUT_TEMPR86[28] , 
        \A_DOUT_TEMPR87[28] , \A_DOUT_TEMPR88[28] , 
        \A_DOUT_TEMPR89[28] , \A_DOUT_TEMPR90[28] , 
        \A_DOUT_TEMPR91[28] , \A_DOUT_TEMPR92[28] , 
        \A_DOUT_TEMPR93[28] , \A_DOUT_TEMPR94[28] , 
        \A_DOUT_TEMPR95[28] , \A_DOUT_TEMPR96[28] , 
        \A_DOUT_TEMPR97[28] , \A_DOUT_TEMPR98[28] , 
        \A_DOUT_TEMPR99[28] , \A_DOUT_TEMPR100[28] , 
        \A_DOUT_TEMPR101[28] , \A_DOUT_TEMPR102[28] , 
        \A_DOUT_TEMPR103[28] , \A_DOUT_TEMPR104[28] , 
        \A_DOUT_TEMPR105[28] , \A_DOUT_TEMPR106[28] , 
        \A_DOUT_TEMPR107[28] , \A_DOUT_TEMPR108[28] , 
        \A_DOUT_TEMPR109[28] , \A_DOUT_TEMPR110[28] , 
        \A_DOUT_TEMPR111[28] , \A_DOUT_TEMPR112[28] , 
        \A_DOUT_TEMPR113[28] , \A_DOUT_TEMPR114[28] , 
        \A_DOUT_TEMPR115[28] , \A_DOUT_TEMPR116[28] , 
        \A_DOUT_TEMPR117[28] , \A_DOUT_TEMPR118[28] , 
        \A_DOUT_TEMPR0[29] , \A_DOUT_TEMPR1[29] , \A_DOUT_TEMPR2[29] , 
        \A_DOUT_TEMPR3[29] , \A_DOUT_TEMPR4[29] , \A_DOUT_TEMPR5[29] , 
        \A_DOUT_TEMPR6[29] , \A_DOUT_TEMPR7[29] , \A_DOUT_TEMPR8[29] , 
        \A_DOUT_TEMPR9[29] , \A_DOUT_TEMPR10[29] , 
        \A_DOUT_TEMPR11[29] , \A_DOUT_TEMPR12[29] , 
        \A_DOUT_TEMPR13[29] , \A_DOUT_TEMPR14[29] , 
        \A_DOUT_TEMPR15[29] , \A_DOUT_TEMPR16[29] , 
        \A_DOUT_TEMPR17[29] , \A_DOUT_TEMPR18[29] , 
        \A_DOUT_TEMPR19[29] , \A_DOUT_TEMPR20[29] , 
        \A_DOUT_TEMPR21[29] , \A_DOUT_TEMPR22[29] , 
        \A_DOUT_TEMPR23[29] , \A_DOUT_TEMPR24[29] , 
        \A_DOUT_TEMPR25[29] , \A_DOUT_TEMPR26[29] , 
        \A_DOUT_TEMPR27[29] , \A_DOUT_TEMPR28[29] , 
        \A_DOUT_TEMPR29[29] , \A_DOUT_TEMPR30[29] , 
        \A_DOUT_TEMPR31[29] , \A_DOUT_TEMPR32[29] , 
        \A_DOUT_TEMPR33[29] , \A_DOUT_TEMPR34[29] , 
        \A_DOUT_TEMPR35[29] , \A_DOUT_TEMPR36[29] , 
        \A_DOUT_TEMPR37[29] , \A_DOUT_TEMPR38[29] , 
        \A_DOUT_TEMPR39[29] , \A_DOUT_TEMPR40[29] , 
        \A_DOUT_TEMPR41[29] , \A_DOUT_TEMPR42[29] , 
        \A_DOUT_TEMPR43[29] , \A_DOUT_TEMPR44[29] , 
        \A_DOUT_TEMPR45[29] , \A_DOUT_TEMPR46[29] , 
        \A_DOUT_TEMPR47[29] , \A_DOUT_TEMPR48[29] , 
        \A_DOUT_TEMPR49[29] , \A_DOUT_TEMPR50[29] , 
        \A_DOUT_TEMPR51[29] , \A_DOUT_TEMPR52[29] , 
        \A_DOUT_TEMPR53[29] , \A_DOUT_TEMPR54[29] , 
        \A_DOUT_TEMPR55[29] , \A_DOUT_TEMPR56[29] , 
        \A_DOUT_TEMPR57[29] , \A_DOUT_TEMPR58[29] , 
        \A_DOUT_TEMPR59[29] , \A_DOUT_TEMPR60[29] , 
        \A_DOUT_TEMPR61[29] , \A_DOUT_TEMPR62[29] , 
        \A_DOUT_TEMPR63[29] , \A_DOUT_TEMPR64[29] , 
        \A_DOUT_TEMPR65[29] , \A_DOUT_TEMPR66[29] , 
        \A_DOUT_TEMPR67[29] , \A_DOUT_TEMPR68[29] , 
        \A_DOUT_TEMPR69[29] , \A_DOUT_TEMPR70[29] , 
        \A_DOUT_TEMPR71[29] , \A_DOUT_TEMPR72[29] , 
        \A_DOUT_TEMPR73[29] , \A_DOUT_TEMPR74[29] , 
        \A_DOUT_TEMPR75[29] , \A_DOUT_TEMPR76[29] , 
        \A_DOUT_TEMPR77[29] , \A_DOUT_TEMPR78[29] , 
        \A_DOUT_TEMPR79[29] , \A_DOUT_TEMPR80[29] , 
        \A_DOUT_TEMPR81[29] , \A_DOUT_TEMPR82[29] , 
        \A_DOUT_TEMPR83[29] , \A_DOUT_TEMPR84[29] , 
        \A_DOUT_TEMPR85[29] , \A_DOUT_TEMPR86[29] , 
        \A_DOUT_TEMPR87[29] , \A_DOUT_TEMPR88[29] , 
        \A_DOUT_TEMPR89[29] , \A_DOUT_TEMPR90[29] , 
        \A_DOUT_TEMPR91[29] , \A_DOUT_TEMPR92[29] , 
        \A_DOUT_TEMPR93[29] , \A_DOUT_TEMPR94[29] , 
        \A_DOUT_TEMPR95[29] , \A_DOUT_TEMPR96[29] , 
        \A_DOUT_TEMPR97[29] , \A_DOUT_TEMPR98[29] , 
        \A_DOUT_TEMPR99[29] , \A_DOUT_TEMPR100[29] , 
        \A_DOUT_TEMPR101[29] , \A_DOUT_TEMPR102[29] , 
        \A_DOUT_TEMPR103[29] , \A_DOUT_TEMPR104[29] , 
        \A_DOUT_TEMPR105[29] , \A_DOUT_TEMPR106[29] , 
        \A_DOUT_TEMPR107[29] , \A_DOUT_TEMPR108[29] , 
        \A_DOUT_TEMPR109[29] , \A_DOUT_TEMPR110[29] , 
        \A_DOUT_TEMPR111[29] , \A_DOUT_TEMPR112[29] , 
        \A_DOUT_TEMPR113[29] , \A_DOUT_TEMPR114[29] , 
        \A_DOUT_TEMPR115[29] , \A_DOUT_TEMPR116[29] , 
        \A_DOUT_TEMPR117[29] , \A_DOUT_TEMPR118[29] , 
        \A_DOUT_TEMPR0[30] , \A_DOUT_TEMPR1[30] , \A_DOUT_TEMPR2[30] , 
        \A_DOUT_TEMPR3[30] , \A_DOUT_TEMPR4[30] , \A_DOUT_TEMPR5[30] , 
        \A_DOUT_TEMPR6[30] , \A_DOUT_TEMPR7[30] , \A_DOUT_TEMPR8[30] , 
        \A_DOUT_TEMPR9[30] , \A_DOUT_TEMPR10[30] , 
        \A_DOUT_TEMPR11[30] , \A_DOUT_TEMPR12[30] , 
        \A_DOUT_TEMPR13[30] , \A_DOUT_TEMPR14[30] , 
        \A_DOUT_TEMPR15[30] , \A_DOUT_TEMPR16[30] , 
        \A_DOUT_TEMPR17[30] , \A_DOUT_TEMPR18[30] , 
        \A_DOUT_TEMPR19[30] , \A_DOUT_TEMPR20[30] , 
        \A_DOUT_TEMPR21[30] , \A_DOUT_TEMPR22[30] , 
        \A_DOUT_TEMPR23[30] , \A_DOUT_TEMPR24[30] , 
        \A_DOUT_TEMPR25[30] , \A_DOUT_TEMPR26[30] , 
        \A_DOUT_TEMPR27[30] , \A_DOUT_TEMPR28[30] , 
        \A_DOUT_TEMPR29[30] , \A_DOUT_TEMPR30[30] , 
        \A_DOUT_TEMPR31[30] , \A_DOUT_TEMPR32[30] , 
        \A_DOUT_TEMPR33[30] , \A_DOUT_TEMPR34[30] , 
        \A_DOUT_TEMPR35[30] , \A_DOUT_TEMPR36[30] , 
        \A_DOUT_TEMPR37[30] , \A_DOUT_TEMPR38[30] , 
        \A_DOUT_TEMPR39[30] , \A_DOUT_TEMPR40[30] , 
        \A_DOUT_TEMPR41[30] , \A_DOUT_TEMPR42[30] , 
        \A_DOUT_TEMPR43[30] , \A_DOUT_TEMPR44[30] , 
        \A_DOUT_TEMPR45[30] , \A_DOUT_TEMPR46[30] , 
        \A_DOUT_TEMPR47[30] , \A_DOUT_TEMPR48[30] , 
        \A_DOUT_TEMPR49[30] , \A_DOUT_TEMPR50[30] , 
        \A_DOUT_TEMPR51[30] , \A_DOUT_TEMPR52[30] , 
        \A_DOUT_TEMPR53[30] , \A_DOUT_TEMPR54[30] , 
        \A_DOUT_TEMPR55[30] , \A_DOUT_TEMPR56[30] , 
        \A_DOUT_TEMPR57[30] , \A_DOUT_TEMPR58[30] , 
        \A_DOUT_TEMPR59[30] , \A_DOUT_TEMPR60[30] , 
        \A_DOUT_TEMPR61[30] , \A_DOUT_TEMPR62[30] , 
        \A_DOUT_TEMPR63[30] , \A_DOUT_TEMPR64[30] , 
        \A_DOUT_TEMPR65[30] , \A_DOUT_TEMPR66[30] , 
        \A_DOUT_TEMPR67[30] , \A_DOUT_TEMPR68[30] , 
        \A_DOUT_TEMPR69[30] , \A_DOUT_TEMPR70[30] , 
        \A_DOUT_TEMPR71[30] , \A_DOUT_TEMPR72[30] , 
        \A_DOUT_TEMPR73[30] , \A_DOUT_TEMPR74[30] , 
        \A_DOUT_TEMPR75[30] , \A_DOUT_TEMPR76[30] , 
        \A_DOUT_TEMPR77[30] , \A_DOUT_TEMPR78[30] , 
        \A_DOUT_TEMPR79[30] , \A_DOUT_TEMPR80[30] , 
        \A_DOUT_TEMPR81[30] , \A_DOUT_TEMPR82[30] , 
        \A_DOUT_TEMPR83[30] , \A_DOUT_TEMPR84[30] , 
        \A_DOUT_TEMPR85[30] , \A_DOUT_TEMPR86[30] , 
        \A_DOUT_TEMPR87[30] , \A_DOUT_TEMPR88[30] , 
        \A_DOUT_TEMPR89[30] , \A_DOUT_TEMPR90[30] , 
        \A_DOUT_TEMPR91[30] , \A_DOUT_TEMPR92[30] , 
        \A_DOUT_TEMPR93[30] , \A_DOUT_TEMPR94[30] , 
        \A_DOUT_TEMPR95[30] , \A_DOUT_TEMPR96[30] , 
        \A_DOUT_TEMPR97[30] , \A_DOUT_TEMPR98[30] , 
        \A_DOUT_TEMPR99[30] , \A_DOUT_TEMPR100[30] , 
        \A_DOUT_TEMPR101[30] , \A_DOUT_TEMPR102[30] , 
        \A_DOUT_TEMPR103[30] , \A_DOUT_TEMPR104[30] , 
        \A_DOUT_TEMPR105[30] , \A_DOUT_TEMPR106[30] , 
        \A_DOUT_TEMPR107[30] , \A_DOUT_TEMPR108[30] , 
        \A_DOUT_TEMPR109[30] , \A_DOUT_TEMPR110[30] , 
        \A_DOUT_TEMPR111[30] , \A_DOUT_TEMPR112[30] , 
        \A_DOUT_TEMPR113[30] , \A_DOUT_TEMPR114[30] , 
        \A_DOUT_TEMPR115[30] , \A_DOUT_TEMPR116[30] , 
        \A_DOUT_TEMPR117[30] , \A_DOUT_TEMPR118[30] , 
        \A_DOUT_TEMPR0[31] , \A_DOUT_TEMPR1[31] , \A_DOUT_TEMPR2[31] , 
        \A_DOUT_TEMPR3[31] , \A_DOUT_TEMPR4[31] , \A_DOUT_TEMPR5[31] , 
        \A_DOUT_TEMPR6[31] , \A_DOUT_TEMPR7[31] , \A_DOUT_TEMPR8[31] , 
        \A_DOUT_TEMPR9[31] , \A_DOUT_TEMPR10[31] , 
        \A_DOUT_TEMPR11[31] , \A_DOUT_TEMPR12[31] , 
        \A_DOUT_TEMPR13[31] , \A_DOUT_TEMPR14[31] , 
        \A_DOUT_TEMPR15[31] , \A_DOUT_TEMPR16[31] , 
        \A_DOUT_TEMPR17[31] , \A_DOUT_TEMPR18[31] , 
        \A_DOUT_TEMPR19[31] , \A_DOUT_TEMPR20[31] , 
        \A_DOUT_TEMPR21[31] , \A_DOUT_TEMPR22[31] , 
        \A_DOUT_TEMPR23[31] , \A_DOUT_TEMPR24[31] , 
        \A_DOUT_TEMPR25[31] , \A_DOUT_TEMPR26[31] , 
        \A_DOUT_TEMPR27[31] , \A_DOUT_TEMPR28[31] , 
        \A_DOUT_TEMPR29[31] , \A_DOUT_TEMPR30[31] , 
        \A_DOUT_TEMPR31[31] , \A_DOUT_TEMPR32[31] , 
        \A_DOUT_TEMPR33[31] , \A_DOUT_TEMPR34[31] , 
        \A_DOUT_TEMPR35[31] , \A_DOUT_TEMPR36[31] , 
        \A_DOUT_TEMPR37[31] , \A_DOUT_TEMPR38[31] , 
        \A_DOUT_TEMPR39[31] , \A_DOUT_TEMPR40[31] , 
        \A_DOUT_TEMPR41[31] , \A_DOUT_TEMPR42[31] , 
        \A_DOUT_TEMPR43[31] , \A_DOUT_TEMPR44[31] , 
        \A_DOUT_TEMPR45[31] , \A_DOUT_TEMPR46[31] , 
        \A_DOUT_TEMPR47[31] , \A_DOUT_TEMPR48[31] , 
        \A_DOUT_TEMPR49[31] , \A_DOUT_TEMPR50[31] , 
        \A_DOUT_TEMPR51[31] , \A_DOUT_TEMPR52[31] , 
        \A_DOUT_TEMPR53[31] , \A_DOUT_TEMPR54[31] , 
        \A_DOUT_TEMPR55[31] , \A_DOUT_TEMPR56[31] , 
        \A_DOUT_TEMPR57[31] , \A_DOUT_TEMPR58[31] , 
        \A_DOUT_TEMPR59[31] , \A_DOUT_TEMPR60[31] , 
        \A_DOUT_TEMPR61[31] , \A_DOUT_TEMPR62[31] , 
        \A_DOUT_TEMPR63[31] , \A_DOUT_TEMPR64[31] , 
        \A_DOUT_TEMPR65[31] , \A_DOUT_TEMPR66[31] , 
        \A_DOUT_TEMPR67[31] , \A_DOUT_TEMPR68[31] , 
        \A_DOUT_TEMPR69[31] , \A_DOUT_TEMPR70[31] , 
        \A_DOUT_TEMPR71[31] , \A_DOUT_TEMPR72[31] , 
        \A_DOUT_TEMPR73[31] , \A_DOUT_TEMPR74[31] , 
        \A_DOUT_TEMPR75[31] , \A_DOUT_TEMPR76[31] , 
        \A_DOUT_TEMPR77[31] , \A_DOUT_TEMPR78[31] , 
        \A_DOUT_TEMPR79[31] , \A_DOUT_TEMPR80[31] , 
        \A_DOUT_TEMPR81[31] , \A_DOUT_TEMPR82[31] , 
        \A_DOUT_TEMPR83[31] , \A_DOUT_TEMPR84[31] , 
        \A_DOUT_TEMPR85[31] , \A_DOUT_TEMPR86[31] , 
        \A_DOUT_TEMPR87[31] , \A_DOUT_TEMPR88[31] , 
        \A_DOUT_TEMPR89[31] , \A_DOUT_TEMPR90[31] , 
        \A_DOUT_TEMPR91[31] , \A_DOUT_TEMPR92[31] , 
        \A_DOUT_TEMPR93[31] , \A_DOUT_TEMPR94[31] , 
        \A_DOUT_TEMPR95[31] , \A_DOUT_TEMPR96[31] , 
        \A_DOUT_TEMPR97[31] , \A_DOUT_TEMPR98[31] , 
        \A_DOUT_TEMPR99[31] , \A_DOUT_TEMPR100[31] , 
        \A_DOUT_TEMPR101[31] , \A_DOUT_TEMPR102[31] , 
        \A_DOUT_TEMPR103[31] , \A_DOUT_TEMPR104[31] , 
        \A_DOUT_TEMPR105[31] , \A_DOUT_TEMPR106[31] , 
        \A_DOUT_TEMPR107[31] , \A_DOUT_TEMPR108[31] , 
        \A_DOUT_TEMPR109[31] , \A_DOUT_TEMPR110[31] , 
        \A_DOUT_TEMPR111[31] , \A_DOUT_TEMPR112[31] , 
        \A_DOUT_TEMPR113[31] , \A_DOUT_TEMPR114[31] , 
        \A_DOUT_TEMPR115[31] , \A_DOUT_TEMPR116[31] , 
        \A_DOUT_TEMPR117[31] , \A_DOUT_TEMPR118[31] , 
        \A_DOUT_TEMPR0[32] , \A_DOUT_TEMPR1[32] , \A_DOUT_TEMPR2[32] , 
        \A_DOUT_TEMPR3[32] , \A_DOUT_TEMPR4[32] , \A_DOUT_TEMPR5[32] , 
        \A_DOUT_TEMPR6[32] , \A_DOUT_TEMPR7[32] , \A_DOUT_TEMPR8[32] , 
        \A_DOUT_TEMPR9[32] , \A_DOUT_TEMPR10[32] , 
        \A_DOUT_TEMPR11[32] , \A_DOUT_TEMPR12[32] , 
        \A_DOUT_TEMPR13[32] , \A_DOUT_TEMPR14[32] , 
        \A_DOUT_TEMPR15[32] , \A_DOUT_TEMPR16[32] , 
        \A_DOUT_TEMPR17[32] , \A_DOUT_TEMPR18[32] , 
        \A_DOUT_TEMPR19[32] , \A_DOUT_TEMPR20[32] , 
        \A_DOUT_TEMPR21[32] , \A_DOUT_TEMPR22[32] , 
        \A_DOUT_TEMPR23[32] , \A_DOUT_TEMPR24[32] , 
        \A_DOUT_TEMPR25[32] , \A_DOUT_TEMPR26[32] , 
        \A_DOUT_TEMPR27[32] , \A_DOUT_TEMPR28[32] , 
        \A_DOUT_TEMPR29[32] , \A_DOUT_TEMPR30[32] , 
        \A_DOUT_TEMPR31[32] , \A_DOUT_TEMPR32[32] , 
        \A_DOUT_TEMPR33[32] , \A_DOUT_TEMPR34[32] , 
        \A_DOUT_TEMPR35[32] , \A_DOUT_TEMPR36[32] , 
        \A_DOUT_TEMPR37[32] , \A_DOUT_TEMPR38[32] , 
        \A_DOUT_TEMPR39[32] , \A_DOUT_TEMPR40[32] , 
        \A_DOUT_TEMPR41[32] , \A_DOUT_TEMPR42[32] , 
        \A_DOUT_TEMPR43[32] , \A_DOUT_TEMPR44[32] , 
        \A_DOUT_TEMPR45[32] , \A_DOUT_TEMPR46[32] , 
        \A_DOUT_TEMPR47[32] , \A_DOUT_TEMPR48[32] , 
        \A_DOUT_TEMPR49[32] , \A_DOUT_TEMPR50[32] , 
        \A_DOUT_TEMPR51[32] , \A_DOUT_TEMPR52[32] , 
        \A_DOUT_TEMPR53[32] , \A_DOUT_TEMPR54[32] , 
        \A_DOUT_TEMPR55[32] , \A_DOUT_TEMPR56[32] , 
        \A_DOUT_TEMPR57[32] , \A_DOUT_TEMPR58[32] , 
        \A_DOUT_TEMPR59[32] , \A_DOUT_TEMPR60[32] , 
        \A_DOUT_TEMPR61[32] , \A_DOUT_TEMPR62[32] , 
        \A_DOUT_TEMPR63[32] , \A_DOUT_TEMPR64[32] , 
        \A_DOUT_TEMPR65[32] , \A_DOUT_TEMPR66[32] , 
        \A_DOUT_TEMPR67[32] , \A_DOUT_TEMPR68[32] , 
        \A_DOUT_TEMPR69[32] , \A_DOUT_TEMPR70[32] , 
        \A_DOUT_TEMPR71[32] , \A_DOUT_TEMPR72[32] , 
        \A_DOUT_TEMPR73[32] , \A_DOUT_TEMPR74[32] , 
        \A_DOUT_TEMPR75[32] , \A_DOUT_TEMPR76[32] , 
        \A_DOUT_TEMPR77[32] , \A_DOUT_TEMPR78[32] , 
        \A_DOUT_TEMPR79[32] , \A_DOUT_TEMPR80[32] , 
        \A_DOUT_TEMPR81[32] , \A_DOUT_TEMPR82[32] , 
        \A_DOUT_TEMPR83[32] , \A_DOUT_TEMPR84[32] , 
        \A_DOUT_TEMPR85[32] , \A_DOUT_TEMPR86[32] , 
        \A_DOUT_TEMPR87[32] , \A_DOUT_TEMPR88[32] , 
        \A_DOUT_TEMPR89[32] , \A_DOUT_TEMPR90[32] , 
        \A_DOUT_TEMPR91[32] , \A_DOUT_TEMPR92[32] , 
        \A_DOUT_TEMPR93[32] , \A_DOUT_TEMPR94[32] , 
        \A_DOUT_TEMPR95[32] , \A_DOUT_TEMPR96[32] , 
        \A_DOUT_TEMPR97[32] , \A_DOUT_TEMPR98[32] , 
        \A_DOUT_TEMPR99[32] , \A_DOUT_TEMPR100[32] , 
        \A_DOUT_TEMPR101[32] , \A_DOUT_TEMPR102[32] , 
        \A_DOUT_TEMPR103[32] , \A_DOUT_TEMPR104[32] , 
        \A_DOUT_TEMPR105[32] , \A_DOUT_TEMPR106[32] , 
        \A_DOUT_TEMPR107[32] , \A_DOUT_TEMPR108[32] , 
        \A_DOUT_TEMPR109[32] , \A_DOUT_TEMPR110[32] , 
        \A_DOUT_TEMPR111[32] , \A_DOUT_TEMPR112[32] , 
        \A_DOUT_TEMPR113[32] , \A_DOUT_TEMPR114[32] , 
        \A_DOUT_TEMPR115[32] , \A_DOUT_TEMPR116[32] , 
        \A_DOUT_TEMPR117[32] , \A_DOUT_TEMPR118[32] , 
        \A_DOUT_TEMPR0[33] , \A_DOUT_TEMPR1[33] , \A_DOUT_TEMPR2[33] , 
        \A_DOUT_TEMPR3[33] , \A_DOUT_TEMPR4[33] , \A_DOUT_TEMPR5[33] , 
        \A_DOUT_TEMPR6[33] , \A_DOUT_TEMPR7[33] , \A_DOUT_TEMPR8[33] , 
        \A_DOUT_TEMPR9[33] , \A_DOUT_TEMPR10[33] , 
        \A_DOUT_TEMPR11[33] , \A_DOUT_TEMPR12[33] , 
        \A_DOUT_TEMPR13[33] , \A_DOUT_TEMPR14[33] , 
        \A_DOUT_TEMPR15[33] , \A_DOUT_TEMPR16[33] , 
        \A_DOUT_TEMPR17[33] , \A_DOUT_TEMPR18[33] , 
        \A_DOUT_TEMPR19[33] , \A_DOUT_TEMPR20[33] , 
        \A_DOUT_TEMPR21[33] , \A_DOUT_TEMPR22[33] , 
        \A_DOUT_TEMPR23[33] , \A_DOUT_TEMPR24[33] , 
        \A_DOUT_TEMPR25[33] , \A_DOUT_TEMPR26[33] , 
        \A_DOUT_TEMPR27[33] , \A_DOUT_TEMPR28[33] , 
        \A_DOUT_TEMPR29[33] , \A_DOUT_TEMPR30[33] , 
        \A_DOUT_TEMPR31[33] , \A_DOUT_TEMPR32[33] , 
        \A_DOUT_TEMPR33[33] , \A_DOUT_TEMPR34[33] , 
        \A_DOUT_TEMPR35[33] , \A_DOUT_TEMPR36[33] , 
        \A_DOUT_TEMPR37[33] , \A_DOUT_TEMPR38[33] , 
        \A_DOUT_TEMPR39[33] , \A_DOUT_TEMPR40[33] , 
        \A_DOUT_TEMPR41[33] , \A_DOUT_TEMPR42[33] , 
        \A_DOUT_TEMPR43[33] , \A_DOUT_TEMPR44[33] , 
        \A_DOUT_TEMPR45[33] , \A_DOUT_TEMPR46[33] , 
        \A_DOUT_TEMPR47[33] , \A_DOUT_TEMPR48[33] , 
        \A_DOUT_TEMPR49[33] , \A_DOUT_TEMPR50[33] , 
        \A_DOUT_TEMPR51[33] , \A_DOUT_TEMPR52[33] , 
        \A_DOUT_TEMPR53[33] , \A_DOUT_TEMPR54[33] , 
        \A_DOUT_TEMPR55[33] , \A_DOUT_TEMPR56[33] , 
        \A_DOUT_TEMPR57[33] , \A_DOUT_TEMPR58[33] , 
        \A_DOUT_TEMPR59[33] , \A_DOUT_TEMPR60[33] , 
        \A_DOUT_TEMPR61[33] , \A_DOUT_TEMPR62[33] , 
        \A_DOUT_TEMPR63[33] , \A_DOUT_TEMPR64[33] , 
        \A_DOUT_TEMPR65[33] , \A_DOUT_TEMPR66[33] , 
        \A_DOUT_TEMPR67[33] , \A_DOUT_TEMPR68[33] , 
        \A_DOUT_TEMPR69[33] , \A_DOUT_TEMPR70[33] , 
        \A_DOUT_TEMPR71[33] , \A_DOUT_TEMPR72[33] , 
        \A_DOUT_TEMPR73[33] , \A_DOUT_TEMPR74[33] , 
        \A_DOUT_TEMPR75[33] , \A_DOUT_TEMPR76[33] , 
        \A_DOUT_TEMPR77[33] , \A_DOUT_TEMPR78[33] , 
        \A_DOUT_TEMPR79[33] , \A_DOUT_TEMPR80[33] , 
        \A_DOUT_TEMPR81[33] , \A_DOUT_TEMPR82[33] , 
        \A_DOUT_TEMPR83[33] , \A_DOUT_TEMPR84[33] , 
        \A_DOUT_TEMPR85[33] , \A_DOUT_TEMPR86[33] , 
        \A_DOUT_TEMPR87[33] , \A_DOUT_TEMPR88[33] , 
        \A_DOUT_TEMPR89[33] , \A_DOUT_TEMPR90[33] , 
        \A_DOUT_TEMPR91[33] , \A_DOUT_TEMPR92[33] , 
        \A_DOUT_TEMPR93[33] , \A_DOUT_TEMPR94[33] , 
        \A_DOUT_TEMPR95[33] , \A_DOUT_TEMPR96[33] , 
        \A_DOUT_TEMPR97[33] , \A_DOUT_TEMPR98[33] , 
        \A_DOUT_TEMPR99[33] , \A_DOUT_TEMPR100[33] , 
        \A_DOUT_TEMPR101[33] , \A_DOUT_TEMPR102[33] , 
        \A_DOUT_TEMPR103[33] , \A_DOUT_TEMPR104[33] , 
        \A_DOUT_TEMPR105[33] , \A_DOUT_TEMPR106[33] , 
        \A_DOUT_TEMPR107[33] , \A_DOUT_TEMPR108[33] , 
        \A_DOUT_TEMPR109[33] , \A_DOUT_TEMPR110[33] , 
        \A_DOUT_TEMPR111[33] , \A_DOUT_TEMPR112[33] , 
        \A_DOUT_TEMPR113[33] , \A_DOUT_TEMPR114[33] , 
        \A_DOUT_TEMPR115[33] , \A_DOUT_TEMPR116[33] , 
        \A_DOUT_TEMPR117[33] , \A_DOUT_TEMPR118[33] , 
        \A_DOUT_TEMPR0[34] , \A_DOUT_TEMPR1[34] , \A_DOUT_TEMPR2[34] , 
        \A_DOUT_TEMPR3[34] , \A_DOUT_TEMPR4[34] , \A_DOUT_TEMPR5[34] , 
        \A_DOUT_TEMPR6[34] , \A_DOUT_TEMPR7[34] , \A_DOUT_TEMPR8[34] , 
        \A_DOUT_TEMPR9[34] , \A_DOUT_TEMPR10[34] , 
        \A_DOUT_TEMPR11[34] , \A_DOUT_TEMPR12[34] , 
        \A_DOUT_TEMPR13[34] , \A_DOUT_TEMPR14[34] , 
        \A_DOUT_TEMPR15[34] , \A_DOUT_TEMPR16[34] , 
        \A_DOUT_TEMPR17[34] , \A_DOUT_TEMPR18[34] , 
        \A_DOUT_TEMPR19[34] , \A_DOUT_TEMPR20[34] , 
        \A_DOUT_TEMPR21[34] , \A_DOUT_TEMPR22[34] , 
        \A_DOUT_TEMPR23[34] , \A_DOUT_TEMPR24[34] , 
        \A_DOUT_TEMPR25[34] , \A_DOUT_TEMPR26[34] , 
        \A_DOUT_TEMPR27[34] , \A_DOUT_TEMPR28[34] , 
        \A_DOUT_TEMPR29[34] , \A_DOUT_TEMPR30[34] , 
        \A_DOUT_TEMPR31[34] , \A_DOUT_TEMPR32[34] , 
        \A_DOUT_TEMPR33[34] , \A_DOUT_TEMPR34[34] , 
        \A_DOUT_TEMPR35[34] , \A_DOUT_TEMPR36[34] , 
        \A_DOUT_TEMPR37[34] , \A_DOUT_TEMPR38[34] , 
        \A_DOUT_TEMPR39[34] , \A_DOUT_TEMPR40[34] , 
        \A_DOUT_TEMPR41[34] , \A_DOUT_TEMPR42[34] , 
        \A_DOUT_TEMPR43[34] , \A_DOUT_TEMPR44[34] , 
        \A_DOUT_TEMPR45[34] , \A_DOUT_TEMPR46[34] , 
        \A_DOUT_TEMPR47[34] , \A_DOUT_TEMPR48[34] , 
        \A_DOUT_TEMPR49[34] , \A_DOUT_TEMPR50[34] , 
        \A_DOUT_TEMPR51[34] , \A_DOUT_TEMPR52[34] , 
        \A_DOUT_TEMPR53[34] , \A_DOUT_TEMPR54[34] , 
        \A_DOUT_TEMPR55[34] , \A_DOUT_TEMPR56[34] , 
        \A_DOUT_TEMPR57[34] , \A_DOUT_TEMPR58[34] , 
        \A_DOUT_TEMPR59[34] , \A_DOUT_TEMPR60[34] , 
        \A_DOUT_TEMPR61[34] , \A_DOUT_TEMPR62[34] , 
        \A_DOUT_TEMPR63[34] , \A_DOUT_TEMPR64[34] , 
        \A_DOUT_TEMPR65[34] , \A_DOUT_TEMPR66[34] , 
        \A_DOUT_TEMPR67[34] , \A_DOUT_TEMPR68[34] , 
        \A_DOUT_TEMPR69[34] , \A_DOUT_TEMPR70[34] , 
        \A_DOUT_TEMPR71[34] , \A_DOUT_TEMPR72[34] , 
        \A_DOUT_TEMPR73[34] , \A_DOUT_TEMPR74[34] , 
        \A_DOUT_TEMPR75[34] , \A_DOUT_TEMPR76[34] , 
        \A_DOUT_TEMPR77[34] , \A_DOUT_TEMPR78[34] , 
        \A_DOUT_TEMPR79[34] , \A_DOUT_TEMPR80[34] , 
        \A_DOUT_TEMPR81[34] , \A_DOUT_TEMPR82[34] , 
        \A_DOUT_TEMPR83[34] , \A_DOUT_TEMPR84[34] , 
        \A_DOUT_TEMPR85[34] , \A_DOUT_TEMPR86[34] , 
        \A_DOUT_TEMPR87[34] , \A_DOUT_TEMPR88[34] , 
        \A_DOUT_TEMPR89[34] , \A_DOUT_TEMPR90[34] , 
        \A_DOUT_TEMPR91[34] , \A_DOUT_TEMPR92[34] , 
        \A_DOUT_TEMPR93[34] , \A_DOUT_TEMPR94[34] , 
        \A_DOUT_TEMPR95[34] , \A_DOUT_TEMPR96[34] , 
        \A_DOUT_TEMPR97[34] , \A_DOUT_TEMPR98[34] , 
        \A_DOUT_TEMPR99[34] , \A_DOUT_TEMPR100[34] , 
        \A_DOUT_TEMPR101[34] , \A_DOUT_TEMPR102[34] , 
        \A_DOUT_TEMPR103[34] , \A_DOUT_TEMPR104[34] , 
        \A_DOUT_TEMPR105[34] , \A_DOUT_TEMPR106[34] , 
        \A_DOUT_TEMPR107[34] , \A_DOUT_TEMPR108[34] , 
        \A_DOUT_TEMPR109[34] , \A_DOUT_TEMPR110[34] , 
        \A_DOUT_TEMPR111[34] , \A_DOUT_TEMPR112[34] , 
        \A_DOUT_TEMPR113[34] , \A_DOUT_TEMPR114[34] , 
        \A_DOUT_TEMPR115[34] , \A_DOUT_TEMPR116[34] , 
        \A_DOUT_TEMPR117[34] , \A_DOUT_TEMPR118[34] , 
        \A_DOUT_TEMPR0[35] , \A_DOUT_TEMPR1[35] , \A_DOUT_TEMPR2[35] , 
        \A_DOUT_TEMPR3[35] , \A_DOUT_TEMPR4[35] , \A_DOUT_TEMPR5[35] , 
        \A_DOUT_TEMPR6[35] , \A_DOUT_TEMPR7[35] , \A_DOUT_TEMPR8[35] , 
        \A_DOUT_TEMPR9[35] , \A_DOUT_TEMPR10[35] , 
        \A_DOUT_TEMPR11[35] , \A_DOUT_TEMPR12[35] , 
        \A_DOUT_TEMPR13[35] , \A_DOUT_TEMPR14[35] , 
        \A_DOUT_TEMPR15[35] , \A_DOUT_TEMPR16[35] , 
        \A_DOUT_TEMPR17[35] , \A_DOUT_TEMPR18[35] , 
        \A_DOUT_TEMPR19[35] , \A_DOUT_TEMPR20[35] , 
        \A_DOUT_TEMPR21[35] , \A_DOUT_TEMPR22[35] , 
        \A_DOUT_TEMPR23[35] , \A_DOUT_TEMPR24[35] , 
        \A_DOUT_TEMPR25[35] , \A_DOUT_TEMPR26[35] , 
        \A_DOUT_TEMPR27[35] , \A_DOUT_TEMPR28[35] , 
        \A_DOUT_TEMPR29[35] , \A_DOUT_TEMPR30[35] , 
        \A_DOUT_TEMPR31[35] , \A_DOUT_TEMPR32[35] , 
        \A_DOUT_TEMPR33[35] , \A_DOUT_TEMPR34[35] , 
        \A_DOUT_TEMPR35[35] , \A_DOUT_TEMPR36[35] , 
        \A_DOUT_TEMPR37[35] , \A_DOUT_TEMPR38[35] , 
        \A_DOUT_TEMPR39[35] , \A_DOUT_TEMPR40[35] , 
        \A_DOUT_TEMPR41[35] , \A_DOUT_TEMPR42[35] , 
        \A_DOUT_TEMPR43[35] , \A_DOUT_TEMPR44[35] , 
        \A_DOUT_TEMPR45[35] , \A_DOUT_TEMPR46[35] , 
        \A_DOUT_TEMPR47[35] , \A_DOUT_TEMPR48[35] , 
        \A_DOUT_TEMPR49[35] , \A_DOUT_TEMPR50[35] , 
        \A_DOUT_TEMPR51[35] , \A_DOUT_TEMPR52[35] , 
        \A_DOUT_TEMPR53[35] , \A_DOUT_TEMPR54[35] , 
        \A_DOUT_TEMPR55[35] , \A_DOUT_TEMPR56[35] , 
        \A_DOUT_TEMPR57[35] , \A_DOUT_TEMPR58[35] , 
        \A_DOUT_TEMPR59[35] , \A_DOUT_TEMPR60[35] , 
        \A_DOUT_TEMPR61[35] , \A_DOUT_TEMPR62[35] , 
        \A_DOUT_TEMPR63[35] , \A_DOUT_TEMPR64[35] , 
        \A_DOUT_TEMPR65[35] , \A_DOUT_TEMPR66[35] , 
        \A_DOUT_TEMPR67[35] , \A_DOUT_TEMPR68[35] , 
        \A_DOUT_TEMPR69[35] , \A_DOUT_TEMPR70[35] , 
        \A_DOUT_TEMPR71[35] , \A_DOUT_TEMPR72[35] , 
        \A_DOUT_TEMPR73[35] , \A_DOUT_TEMPR74[35] , 
        \A_DOUT_TEMPR75[35] , \A_DOUT_TEMPR76[35] , 
        \A_DOUT_TEMPR77[35] , \A_DOUT_TEMPR78[35] , 
        \A_DOUT_TEMPR79[35] , \A_DOUT_TEMPR80[35] , 
        \A_DOUT_TEMPR81[35] , \A_DOUT_TEMPR82[35] , 
        \A_DOUT_TEMPR83[35] , \A_DOUT_TEMPR84[35] , 
        \A_DOUT_TEMPR85[35] , \A_DOUT_TEMPR86[35] , 
        \A_DOUT_TEMPR87[35] , \A_DOUT_TEMPR88[35] , 
        \A_DOUT_TEMPR89[35] , \A_DOUT_TEMPR90[35] , 
        \A_DOUT_TEMPR91[35] , \A_DOUT_TEMPR92[35] , 
        \A_DOUT_TEMPR93[35] , \A_DOUT_TEMPR94[35] , 
        \A_DOUT_TEMPR95[35] , \A_DOUT_TEMPR96[35] , 
        \A_DOUT_TEMPR97[35] , \A_DOUT_TEMPR98[35] , 
        \A_DOUT_TEMPR99[35] , \A_DOUT_TEMPR100[35] , 
        \A_DOUT_TEMPR101[35] , \A_DOUT_TEMPR102[35] , 
        \A_DOUT_TEMPR103[35] , \A_DOUT_TEMPR104[35] , 
        \A_DOUT_TEMPR105[35] , \A_DOUT_TEMPR106[35] , 
        \A_DOUT_TEMPR107[35] , \A_DOUT_TEMPR108[35] , 
        \A_DOUT_TEMPR109[35] , \A_DOUT_TEMPR110[35] , 
        \A_DOUT_TEMPR111[35] , \A_DOUT_TEMPR112[35] , 
        \A_DOUT_TEMPR113[35] , \A_DOUT_TEMPR114[35] , 
        \A_DOUT_TEMPR115[35] , \A_DOUT_TEMPR116[35] , 
        \A_DOUT_TEMPR117[35] , \A_DOUT_TEMPR118[35] , 
        \A_DOUT_TEMPR0[36] , \A_DOUT_TEMPR1[36] , \A_DOUT_TEMPR2[36] , 
        \A_DOUT_TEMPR3[36] , \A_DOUT_TEMPR4[36] , \A_DOUT_TEMPR5[36] , 
        \A_DOUT_TEMPR6[36] , \A_DOUT_TEMPR7[36] , \A_DOUT_TEMPR8[36] , 
        \A_DOUT_TEMPR9[36] , \A_DOUT_TEMPR10[36] , 
        \A_DOUT_TEMPR11[36] , \A_DOUT_TEMPR12[36] , 
        \A_DOUT_TEMPR13[36] , \A_DOUT_TEMPR14[36] , 
        \A_DOUT_TEMPR15[36] , \A_DOUT_TEMPR16[36] , 
        \A_DOUT_TEMPR17[36] , \A_DOUT_TEMPR18[36] , 
        \A_DOUT_TEMPR19[36] , \A_DOUT_TEMPR20[36] , 
        \A_DOUT_TEMPR21[36] , \A_DOUT_TEMPR22[36] , 
        \A_DOUT_TEMPR23[36] , \A_DOUT_TEMPR24[36] , 
        \A_DOUT_TEMPR25[36] , \A_DOUT_TEMPR26[36] , 
        \A_DOUT_TEMPR27[36] , \A_DOUT_TEMPR28[36] , 
        \A_DOUT_TEMPR29[36] , \A_DOUT_TEMPR30[36] , 
        \A_DOUT_TEMPR31[36] , \A_DOUT_TEMPR32[36] , 
        \A_DOUT_TEMPR33[36] , \A_DOUT_TEMPR34[36] , 
        \A_DOUT_TEMPR35[36] , \A_DOUT_TEMPR36[36] , 
        \A_DOUT_TEMPR37[36] , \A_DOUT_TEMPR38[36] , 
        \A_DOUT_TEMPR39[36] , \A_DOUT_TEMPR40[36] , 
        \A_DOUT_TEMPR41[36] , \A_DOUT_TEMPR42[36] , 
        \A_DOUT_TEMPR43[36] , \A_DOUT_TEMPR44[36] , 
        \A_DOUT_TEMPR45[36] , \A_DOUT_TEMPR46[36] , 
        \A_DOUT_TEMPR47[36] , \A_DOUT_TEMPR48[36] , 
        \A_DOUT_TEMPR49[36] , \A_DOUT_TEMPR50[36] , 
        \A_DOUT_TEMPR51[36] , \A_DOUT_TEMPR52[36] , 
        \A_DOUT_TEMPR53[36] , \A_DOUT_TEMPR54[36] , 
        \A_DOUT_TEMPR55[36] , \A_DOUT_TEMPR56[36] , 
        \A_DOUT_TEMPR57[36] , \A_DOUT_TEMPR58[36] , 
        \A_DOUT_TEMPR59[36] , \A_DOUT_TEMPR60[36] , 
        \A_DOUT_TEMPR61[36] , \A_DOUT_TEMPR62[36] , 
        \A_DOUT_TEMPR63[36] , \A_DOUT_TEMPR64[36] , 
        \A_DOUT_TEMPR65[36] , \A_DOUT_TEMPR66[36] , 
        \A_DOUT_TEMPR67[36] , \A_DOUT_TEMPR68[36] , 
        \A_DOUT_TEMPR69[36] , \A_DOUT_TEMPR70[36] , 
        \A_DOUT_TEMPR71[36] , \A_DOUT_TEMPR72[36] , 
        \A_DOUT_TEMPR73[36] , \A_DOUT_TEMPR74[36] , 
        \A_DOUT_TEMPR75[36] , \A_DOUT_TEMPR76[36] , 
        \A_DOUT_TEMPR77[36] , \A_DOUT_TEMPR78[36] , 
        \A_DOUT_TEMPR79[36] , \A_DOUT_TEMPR80[36] , 
        \A_DOUT_TEMPR81[36] , \A_DOUT_TEMPR82[36] , 
        \A_DOUT_TEMPR83[36] , \A_DOUT_TEMPR84[36] , 
        \A_DOUT_TEMPR85[36] , \A_DOUT_TEMPR86[36] , 
        \A_DOUT_TEMPR87[36] , \A_DOUT_TEMPR88[36] , 
        \A_DOUT_TEMPR89[36] , \A_DOUT_TEMPR90[36] , 
        \A_DOUT_TEMPR91[36] , \A_DOUT_TEMPR92[36] , 
        \A_DOUT_TEMPR93[36] , \A_DOUT_TEMPR94[36] , 
        \A_DOUT_TEMPR95[36] , \A_DOUT_TEMPR96[36] , 
        \A_DOUT_TEMPR97[36] , \A_DOUT_TEMPR98[36] , 
        \A_DOUT_TEMPR99[36] , \A_DOUT_TEMPR100[36] , 
        \A_DOUT_TEMPR101[36] , \A_DOUT_TEMPR102[36] , 
        \A_DOUT_TEMPR103[36] , \A_DOUT_TEMPR104[36] , 
        \A_DOUT_TEMPR105[36] , \A_DOUT_TEMPR106[36] , 
        \A_DOUT_TEMPR107[36] , \A_DOUT_TEMPR108[36] , 
        \A_DOUT_TEMPR109[36] , \A_DOUT_TEMPR110[36] , 
        \A_DOUT_TEMPR111[36] , \A_DOUT_TEMPR112[36] , 
        \A_DOUT_TEMPR113[36] , \A_DOUT_TEMPR114[36] , 
        \A_DOUT_TEMPR115[36] , \A_DOUT_TEMPR116[36] , 
        \A_DOUT_TEMPR117[36] , \A_DOUT_TEMPR118[36] , 
        \A_DOUT_TEMPR0[37] , \A_DOUT_TEMPR1[37] , \A_DOUT_TEMPR2[37] , 
        \A_DOUT_TEMPR3[37] , \A_DOUT_TEMPR4[37] , \A_DOUT_TEMPR5[37] , 
        \A_DOUT_TEMPR6[37] , \A_DOUT_TEMPR7[37] , \A_DOUT_TEMPR8[37] , 
        \A_DOUT_TEMPR9[37] , \A_DOUT_TEMPR10[37] , 
        \A_DOUT_TEMPR11[37] , \A_DOUT_TEMPR12[37] , 
        \A_DOUT_TEMPR13[37] , \A_DOUT_TEMPR14[37] , 
        \A_DOUT_TEMPR15[37] , \A_DOUT_TEMPR16[37] , 
        \A_DOUT_TEMPR17[37] , \A_DOUT_TEMPR18[37] , 
        \A_DOUT_TEMPR19[37] , \A_DOUT_TEMPR20[37] , 
        \A_DOUT_TEMPR21[37] , \A_DOUT_TEMPR22[37] , 
        \A_DOUT_TEMPR23[37] , \A_DOUT_TEMPR24[37] , 
        \A_DOUT_TEMPR25[37] , \A_DOUT_TEMPR26[37] , 
        \A_DOUT_TEMPR27[37] , \A_DOUT_TEMPR28[37] , 
        \A_DOUT_TEMPR29[37] , \A_DOUT_TEMPR30[37] , 
        \A_DOUT_TEMPR31[37] , \A_DOUT_TEMPR32[37] , 
        \A_DOUT_TEMPR33[37] , \A_DOUT_TEMPR34[37] , 
        \A_DOUT_TEMPR35[37] , \A_DOUT_TEMPR36[37] , 
        \A_DOUT_TEMPR37[37] , \A_DOUT_TEMPR38[37] , 
        \A_DOUT_TEMPR39[37] , \A_DOUT_TEMPR40[37] , 
        \A_DOUT_TEMPR41[37] , \A_DOUT_TEMPR42[37] , 
        \A_DOUT_TEMPR43[37] , \A_DOUT_TEMPR44[37] , 
        \A_DOUT_TEMPR45[37] , \A_DOUT_TEMPR46[37] , 
        \A_DOUT_TEMPR47[37] , \A_DOUT_TEMPR48[37] , 
        \A_DOUT_TEMPR49[37] , \A_DOUT_TEMPR50[37] , 
        \A_DOUT_TEMPR51[37] , \A_DOUT_TEMPR52[37] , 
        \A_DOUT_TEMPR53[37] , \A_DOUT_TEMPR54[37] , 
        \A_DOUT_TEMPR55[37] , \A_DOUT_TEMPR56[37] , 
        \A_DOUT_TEMPR57[37] , \A_DOUT_TEMPR58[37] , 
        \A_DOUT_TEMPR59[37] , \A_DOUT_TEMPR60[37] , 
        \A_DOUT_TEMPR61[37] , \A_DOUT_TEMPR62[37] , 
        \A_DOUT_TEMPR63[37] , \A_DOUT_TEMPR64[37] , 
        \A_DOUT_TEMPR65[37] , \A_DOUT_TEMPR66[37] , 
        \A_DOUT_TEMPR67[37] , \A_DOUT_TEMPR68[37] , 
        \A_DOUT_TEMPR69[37] , \A_DOUT_TEMPR70[37] , 
        \A_DOUT_TEMPR71[37] , \A_DOUT_TEMPR72[37] , 
        \A_DOUT_TEMPR73[37] , \A_DOUT_TEMPR74[37] , 
        \A_DOUT_TEMPR75[37] , \A_DOUT_TEMPR76[37] , 
        \A_DOUT_TEMPR77[37] , \A_DOUT_TEMPR78[37] , 
        \A_DOUT_TEMPR79[37] , \A_DOUT_TEMPR80[37] , 
        \A_DOUT_TEMPR81[37] , \A_DOUT_TEMPR82[37] , 
        \A_DOUT_TEMPR83[37] , \A_DOUT_TEMPR84[37] , 
        \A_DOUT_TEMPR85[37] , \A_DOUT_TEMPR86[37] , 
        \A_DOUT_TEMPR87[37] , \A_DOUT_TEMPR88[37] , 
        \A_DOUT_TEMPR89[37] , \A_DOUT_TEMPR90[37] , 
        \A_DOUT_TEMPR91[37] , \A_DOUT_TEMPR92[37] , 
        \A_DOUT_TEMPR93[37] , \A_DOUT_TEMPR94[37] , 
        \A_DOUT_TEMPR95[37] , \A_DOUT_TEMPR96[37] , 
        \A_DOUT_TEMPR97[37] , \A_DOUT_TEMPR98[37] , 
        \A_DOUT_TEMPR99[37] , \A_DOUT_TEMPR100[37] , 
        \A_DOUT_TEMPR101[37] , \A_DOUT_TEMPR102[37] , 
        \A_DOUT_TEMPR103[37] , \A_DOUT_TEMPR104[37] , 
        \A_DOUT_TEMPR105[37] , \A_DOUT_TEMPR106[37] , 
        \A_DOUT_TEMPR107[37] , \A_DOUT_TEMPR108[37] , 
        \A_DOUT_TEMPR109[37] , \A_DOUT_TEMPR110[37] , 
        \A_DOUT_TEMPR111[37] , \A_DOUT_TEMPR112[37] , 
        \A_DOUT_TEMPR113[37] , \A_DOUT_TEMPR114[37] , 
        \A_DOUT_TEMPR115[37] , \A_DOUT_TEMPR116[37] , 
        \A_DOUT_TEMPR117[37] , \A_DOUT_TEMPR118[37] , 
        \A_DOUT_TEMPR0[38] , \A_DOUT_TEMPR1[38] , \A_DOUT_TEMPR2[38] , 
        \A_DOUT_TEMPR3[38] , \A_DOUT_TEMPR4[38] , \A_DOUT_TEMPR5[38] , 
        \A_DOUT_TEMPR6[38] , \A_DOUT_TEMPR7[38] , \A_DOUT_TEMPR8[38] , 
        \A_DOUT_TEMPR9[38] , \A_DOUT_TEMPR10[38] , 
        \A_DOUT_TEMPR11[38] , \A_DOUT_TEMPR12[38] , 
        \A_DOUT_TEMPR13[38] , \A_DOUT_TEMPR14[38] , 
        \A_DOUT_TEMPR15[38] , \A_DOUT_TEMPR16[38] , 
        \A_DOUT_TEMPR17[38] , \A_DOUT_TEMPR18[38] , 
        \A_DOUT_TEMPR19[38] , \A_DOUT_TEMPR20[38] , 
        \A_DOUT_TEMPR21[38] , \A_DOUT_TEMPR22[38] , 
        \A_DOUT_TEMPR23[38] , \A_DOUT_TEMPR24[38] , 
        \A_DOUT_TEMPR25[38] , \A_DOUT_TEMPR26[38] , 
        \A_DOUT_TEMPR27[38] , \A_DOUT_TEMPR28[38] , 
        \A_DOUT_TEMPR29[38] , \A_DOUT_TEMPR30[38] , 
        \A_DOUT_TEMPR31[38] , \A_DOUT_TEMPR32[38] , 
        \A_DOUT_TEMPR33[38] , \A_DOUT_TEMPR34[38] , 
        \A_DOUT_TEMPR35[38] , \A_DOUT_TEMPR36[38] , 
        \A_DOUT_TEMPR37[38] , \A_DOUT_TEMPR38[38] , 
        \A_DOUT_TEMPR39[38] , \A_DOUT_TEMPR40[38] , 
        \A_DOUT_TEMPR41[38] , \A_DOUT_TEMPR42[38] , 
        \A_DOUT_TEMPR43[38] , \A_DOUT_TEMPR44[38] , 
        \A_DOUT_TEMPR45[38] , \A_DOUT_TEMPR46[38] , 
        \A_DOUT_TEMPR47[38] , \A_DOUT_TEMPR48[38] , 
        \A_DOUT_TEMPR49[38] , \A_DOUT_TEMPR50[38] , 
        \A_DOUT_TEMPR51[38] , \A_DOUT_TEMPR52[38] , 
        \A_DOUT_TEMPR53[38] , \A_DOUT_TEMPR54[38] , 
        \A_DOUT_TEMPR55[38] , \A_DOUT_TEMPR56[38] , 
        \A_DOUT_TEMPR57[38] , \A_DOUT_TEMPR58[38] , 
        \A_DOUT_TEMPR59[38] , \A_DOUT_TEMPR60[38] , 
        \A_DOUT_TEMPR61[38] , \A_DOUT_TEMPR62[38] , 
        \A_DOUT_TEMPR63[38] , \A_DOUT_TEMPR64[38] , 
        \A_DOUT_TEMPR65[38] , \A_DOUT_TEMPR66[38] , 
        \A_DOUT_TEMPR67[38] , \A_DOUT_TEMPR68[38] , 
        \A_DOUT_TEMPR69[38] , \A_DOUT_TEMPR70[38] , 
        \A_DOUT_TEMPR71[38] , \A_DOUT_TEMPR72[38] , 
        \A_DOUT_TEMPR73[38] , \A_DOUT_TEMPR74[38] , 
        \A_DOUT_TEMPR75[38] , \A_DOUT_TEMPR76[38] , 
        \A_DOUT_TEMPR77[38] , \A_DOUT_TEMPR78[38] , 
        \A_DOUT_TEMPR79[38] , \A_DOUT_TEMPR80[38] , 
        \A_DOUT_TEMPR81[38] , \A_DOUT_TEMPR82[38] , 
        \A_DOUT_TEMPR83[38] , \A_DOUT_TEMPR84[38] , 
        \A_DOUT_TEMPR85[38] , \A_DOUT_TEMPR86[38] , 
        \A_DOUT_TEMPR87[38] , \A_DOUT_TEMPR88[38] , 
        \A_DOUT_TEMPR89[38] , \A_DOUT_TEMPR90[38] , 
        \A_DOUT_TEMPR91[38] , \A_DOUT_TEMPR92[38] , 
        \A_DOUT_TEMPR93[38] , \A_DOUT_TEMPR94[38] , 
        \A_DOUT_TEMPR95[38] , \A_DOUT_TEMPR96[38] , 
        \A_DOUT_TEMPR97[38] , \A_DOUT_TEMPR98[38] , 
        \A_DOUT_TEMPR99[38] , \A_DOUT_TEMPR100[38] , 
        \A_DOUT_TEMPR101[38] , \A_DOUT_TEMPR102[38] , 
        \A_DOUT_TEMPR103[38] , \A_DOUT_TEMPR104[38] , 
        \A_DOUT_TEMPR105[38] , \A_DOUT_TEMPR106[38] , 
        \A_DOUT_TEMPR107[38] , \A_DOUT_TEMPR108[38] , 
        \A_DOUT_TEMPR109[38] , \A_DOUT_TEMPR110[38] , 
        \A_DOUT_TEMPR111[38] , \A_DOUT_TEMPR112[38] , 
        \A_DOUT_TEMPR113[38] , \A_DOUT_TEMPR114[38] , 
        \A_DOUT_TEMPR115[38] , \A_DOUT_TEMPR116[38] , 
        \A_DOUT_TEMPR117[38] , \A_DOUT_TEMPR118[38] , 
        \A_DOUT_TEMPR0[39] , \A_DOUT_TEMPR1[39] , \A_DOUT_TEMPR2[39] , 
        \A_DOUT_TEMPR3[39] , \A_DOUT_TEMPR4[39] , \A_DOUT_TEMPR5[39] , 
        \A_DOUT_TEMPR6[39] , \A_DOUT_TEMPR7[39] , \A_DOUT_TEMPR8[39] , 
        \A_DOUT_TEMPR9[39] , \A_DOUT_TEMPR10[39] , 
        \A_DOUT_TEMPR11[39] , \A_DOUT_TEMPR12[39] , 
        \A_DOUT_TEMPR13[39] , \A_DOUT_TEMPR14[39] , 
        \A_DOUT_TEMPR15[39] , \A_DOUT_TEMPR16[39] , 
        \A_DOUT_TEMPR17[39] , \A_DOUT_TEMPR18[39] , 
        \A_DOUT_TEMPR19[39] , \A_DOUT_TEMPR20[39] , 
        \A_DOUT_TEMPR21[39] , \A_DOUT_TEMPR22[39] , 
        \A_DOUT_TEMPR23[39] , \A_DOUT_TEMPR24[39] , 
        \A_DOUT_TEMPR25[39] , \A_DOUT_TEMPR26[39] , 
        \A_DOUT_TEMPR27[39] , \A_DOUT_TEMPR28[39] , 
        \A_DOUT_TEMPR29[39] , \A_DOUT_TEMPR30[39] , 
        \A_DOUT_TEMPR31[39] , \A_DOUT_TEMPR32[39] , 
        \A_DOUT_TEMPR33[39] , \A_DOUT_TEMPR34[39] , 
        \A_DOUT_TEMPR35[39] , \A_DOUT_TEMPR36[39] , 
        \A_DOUT_TEMPR37[39] , \A_DOUT_TEMPR38[39] , 
        \A_DOUT_TEMPR39[39] , \A_DOUT_TEMPR40[39] , 
        \A_DOUT_TEMPR41[39] , \A_DOUT_TEMPR42[39] , 
        \A_DOUT_TEMPR43[39] , \A_DOUT_TEMPR44[39] , 
        \A_DOUT_TEMPR45[39] , \A_DOUT_TEMPR46[39] , 
        \A_DOUT_TEMPR47[39] , \A_DOUT_TEMPR48[39] , 
        \A_DOUT_TEMPR49[39] , \A_DOUT_TEMPR50[39] , 
        \A_DOUT_TEMPR51[39] , \A_DOUT_TEMPR52[39] , 
        \A_DOUT_TEMPR53[39] , \A_DOUT_TEMPR54[39] , 
        \A_DOUT_TEMPR55[39] , \A_DOUT_TEMPR56[39] , 
        \A_DOUT_TEMPR57[39] , \A_DOUT_TEMPR58[39] , 
        \A_DOUT_TEMPR59[39] , \A_DOUT_TEMPR60[39] , 
        \A_DOUT_TEMPR61[39] , \A_DOUT_TEMPR62[39] , 
        \A_DOUT_TEMPR63[39] , \A_DOUT_TEMPR64[39] , 
        \A_DOUT_TEMPR65[39] , \A_DOUT_TEMPR66[39] , 
        \A_DOUT_TEMPR67[39] , \A_DOUT_TEMPR68[39] , 
        \A_DOUT_TEMPR69[39] , \A_DOUT_TEMPR70[39] , 
        \A_DOUT_TEMPR71[39] , \A_DOUT_TEMPR72[39] , 
        \A_DOUT_TEMPR73[39] , \A_DOUT_TEMPR74[39] , 
        \A_DOUT_TEMPR75[39] , \A_DOUT_TEMPR76[39] , 
        \A_DOUT_TEMPR77[39] , \A_DOUT_TEMPR78[39] , 
        \A_DOUT_TEMPR79[39] , \A_DOUT_TEMPR80[39] , 
        \A_DOUT_TEMPR81[39] , \A_DOUT_TEMPR82[39] , 
        \A_DOUT_TEMPR83[39] , \A_DOUT_TEMPR84[39] , 
        \A_DOUT_TEMPR85[39] , \A_DOUT_TEMPR86[39] , 
        \A_DOUT_TEMPR87[39] , \A_DOUT_TEMPR88[39] , 
        \A_DOUT_TEMPR89[39] , \A_DOUT_TEMPR90[39] , 
        \A_DOUT_TEMPR91[39] , \A_DOUT_TEMPR92[39] , 
        \A_DOUT_TEMPR93[39] , \A_DOUT_TEMPR94[39] , 
        \A_DOUT_TEMPR95[39] , \A_DOUT_TEMPR96[39] , 
        \A_DOUT_TEMPR97[39] , \A_DOUT_TEMPR98[39] , 
        \A_DOUT_TEMPR99[39] , \A_DOUT_TEMPR100[39] , 
        \A_DOUT_TEMPR101[39] , \A_DOUT_TEMPR102[39] , 
        \A_DOUT_TEMPR103[39] , \A_DOUT_TEMPR104[39] , 
        \A_DOUT_TEMPR105[39] , \A_DOUT_TEMPR106[39] , 
        \A_DOUT_TEMPR107[39] , \A_DOUT_TEMPR108[39] , 
        \A_DOUT_TEMPR109[39] , \A_DOUT_TEMPR110[39] , 
        \A_DOUT_TEMPR111[39] , \A_DOUT_TEMPR112[39] , 
        \A_DOUT_TEMPR113[39] , \A_DOUT_TEMPR114[39] , 
        \A_DOUT_TEMPR115[39] , \A_DOUT_TEMPR116[39] , 
        \A_DOUT_TEMPR117[39] , \A_DOUT_TEMPR118[39] , \BLKX0[0] , 
        \BLKY0[0] , \BLKX1[0] , \BLKY1[0] , \BLKX2[0] , \BLKX2[1] , 
        \BLKX2[2] , \BLKX2[3] , \BLKX2[4] , \BLKX2[5] , \BLKX2[6] , 
        \BLKX2[7] , \BLKX2[8] , \BLKX2[9] , \BLKX2[10] , \BLKX2[11] , 
        \BLKX2[12] , \BLKX2[13] , \BLKX2[14] , \BLKX2[15] , 
        \BLKX2[16] , \BLKX2[17] , \BLKX2[18] , \BLKX2[19] , 
        \BLKX2[20] , \BLKX2[21] , \BLKX2[22] , \BLKX2[23] , 
        \BLKX2[24] , \BLKX2[25] , \BLKX2[26] , \BLKX2[27] , 
        \BLKX2[28] , \BLKX2[29] , \BLKY2[0] , \BLKY2[1] , \BLKY2[2] , 
        \BLKY2[3] , \BLKY2[4] , \BLKY2[5] , \BLKY2[6] , \BLKY2[7] , 
        \BLKY2[8] , \BLKY2[9] , \BLKY2[10] , \BLKY2[11] , \BLKY2[12] , 
        \BLKY2[13] , \BLKY2[14] , \BLKY2[15] , \BLKY2[16] , 
        \BLKY2[17] , \BLKY2[18] , \BLKY2[19] , \BLKY2[20] , 
        \BLKY2[21] , \BLKY2[22] , \BLKY2[23] , \BLKY2[24] , 
        \BLKY2[25] , \BLKY2[26] , \BLKY2[27] , \BLKY2[28] , 
        \BLKY2[29] , \ACCESS_BUSY[0][0] , \ACCESS_BUSY[0][1] , 
        \ACCESS_BUSY[0][2] , \ACCESS_BUSY[0][3] , \ACCESS_BUSY[0][4] , 
        \ACCESS_BUSY[0][5] , \ACCESS_BUSY[0][6] , \ACCESS_BUSY[0][7] , 
        \ACCESS_BUSY[1][0] , \ACCESS_BUSY[1][1] , \ACCESS_BUSY[1][2] , 
        \ACCESS_BUSY[1][3] , \ACCESS_BUSY[1][4] , \ACCESS_BUSY[1][5] , 
        \ACCESS_BUSY[1][6] , \ACCESS_BUSY[1][7] , \ACCESS_BUSY[2][0] , 
        \ACCESS_BUSY[2][1] , \ACCESS_BUSY[2][2] , \ACCESS_BUSY[2][3] , 
        \ACCESS_BUSY[2][4] , \ACCESS_BUSY[2][5] , \ACCESS_BUSY[2][6] , 
        \ACCESS_BUSY[2][7] , \ACCESS_BUSY[3][0] , \ACCESS_BUSY[3][1] , 
        \ACCESS_BUSY[3][2] , \ACCESS_BUSY[3][3] , \ACCESS_BUSY[3][4] , 
        \ACCESS_BUSY[3][5] , \ACCESS_BUSY[3][6] , \ACCESS_BUSY[3][7] , 
        \ACCESS_BUSY[4][0] , \ACCESS_BUSY[4][1] , \ACCESS_BUSY[4][2] , 
        \ACCESS_BUSY[4][3] , \ACCESS_BUSY[4][4] , \ACCESS_BUSY[4][5] , 
        \ACCESS_BUSY[4][6] , \ACCESS_BUSY[4][7] , \ACCESS_BUSY[5][0] , 
        \ACCESS_BUSY[5][1] , \ACCESS_BUSY[5][2] , \ACCESS_BUSY[5][3] , 
        \ACCESS_BUSY[5][4] , \ACCESS_BUSY[5][5] , \ACCESS_BUSY[5][6] , 
        \ACCESS_BUSY[5][7] , \ACCESS_BUSY[6][0] , \ACCESS_BUSY[6][1] , 
        \ACCESS_BUSY[6][2] , \ACCESS_BUSY[6][3] , \ACCESS_BUSY[6][4] , 
        \ACCESS_BUSY[6][5] , \ACCESS_BUSY[6][6] , \ACCESS_BUSY[6][7] , 
        \ACCESS_BUSY[7][0] , \ACCESS_BUSY[7][1] , \ACCESS_BUSY[7][2] , 
        \ACCESS_BUSY[7][3] , \ACCESS_BUSY[7][4] , \ACCESS_BUSY[7][5] , 
        \ACCESS_BUSY[7][6] , \ACCESS_BUSY[7][7] , \ACCESS_BUSY[8][0] , 
        \ACCESS_BUSY[8][1] , \ACCESS_BUSY[8][2] , \ACCESS_BUSY[8][3] , 
        \ACCESS_BUSY[8][4] , \ACCESS_BUSY[8][5] , \ACCESS_BUSY[8][6] , 
        \ACCESS_BUSY[8][7] , \ACCESS_BUSY[9][0] , \ACCESS_BUSY[9][1] , 
        \ACCESS_BUSY[9][2] , \ACCESS_BUSY[9][3] , \ACCESS_BUSY[9][4] , 
        \ACCESS_BUSY[9][5] , \ACCESS_BUSY[9][6] , \ACCESS_BUSY[9][7] , 
        \ACCESS_BUSY[10][0] , \ACCESS_BUSY[10][1] , 
        \ACCESS_BUSY[10][2] , \ACCESS_BUSY[10][3] , 
        \ACCESS_BUSY[10][4] , \ACCESS_BUSY[10][5] , 
        \ACCESS_BUSY[10][6] , \ACCESS_BUSY[10][7] , 
        \ACCESS_BUSY[11][0] , \ACCESS_BUSY[11][1] , 
        \ACCESS_BUSY[11][2] , \ACCESS_BUSY[11][3] , 
        \ACCESS_BUSY[11][4] , \ACCESS_BUSY[11][5] , 
        \ACCESS_BUSY[11][6] , \ACCESS_BUSY[11][7] , 
        \ACCESS_BUSY[12][0] , \ACCESS_BUSY[12][1] , 
        \ACCESS_BUSY[12][2] , \ACCESS_BUSY[12][3] , 
        \ACCESS_BUSY[12][4] , \ACCESS_BUSY[12][5] , 
        \ACCESS_BUSY[12][6] , \ACCESS_BUSY[12][7] , 
        \ACCESS_BUSY[13][0] , \ACCESS_BUSY[13][1] , 
        \ACCESS_BUSY[13][2] , \ACCESS_BUSY[13][3] , 
        \ACCESS_BUSY[13][4] , \ACCESS_BUSY[13][5] , 
        \ACCESS_BUSY[13][6] , \ACCESS_BUSY[13][7] , 
        \ACCESS_BUSY[14][0] , \ACCESS_BUSY[14][1] , 
        \ACCESS_BUSY[14][2] , \ACCESS_BUSY[14][3] , 
        \ACCESS_BUSY[14][4] , \ACCESS_BUSY[14][5] , 
        \ACCESS_BUSY[14][6] , \ACCESS_BUSY[14][7] , 
        \ACCESS_BUSY[15][0] , \ACCESS_BUSY[15][1] , 
        \ACCESS_BUSY[15][2] , \ACCESS_BUSY[15][3] , 
        \ACCESS_BUSY[15][4] , \ACCESS_BUSY[15][5] , 
        \ACCESS_BUSY[15][6] , \ACCESS_BUSY[15][7] , 
        \ACCESS_BUSY[16][0] , \ACCESS_BUSY[16][1] , 
        \ACCESS_BUSY[16][2] , \ACCESS_BUSY[16][3] , 
        \ACCESS_BUSY[16][4] , \ACCESS_BUSY[16][5] , 
        \ACCESS_BUSY[16][6] , \ACCESS_BUSY[16][7] , 
        \ACCESS_BUSY[17][0] , \ACCESS_BUSY[17][1] , 
        \ACCESS_BUSY[17][2] , \ACCESS_BUSY[17][3] , 
        \ACCESS_BUSY[17][4] , \ACCESS_BUSY[17][5] , 
        \ACCESS_BUSY[17][6] , \ACCESS_BUSY[17][7] , 
        \ACCESS_BUSY[18][0] , \ACCESS_BUSY[18][1] , 
        \ACCESS_BUSY[18][2] , \ACCESS_BUSY[18][3] , 
        \ACCESS_BUSY[18][4] , \ACCESS_BUSY[18][5] , 
        \ACCESS_BUSY[18][6] , \ACCESS_BUSY[18][7] , 
        \ACCESS_BUSY[19][0] , \ACCESS_BUSY[19][1] , 
        \ACCESS_BUSY[19][2] , \ACCESS_BUSY[19][3] , 
        \ACCESS_BUSY[19][4] , \ACCESS_BUSY[19][5] , 
        \ACCESS_BUSY[19][6] , \ACCESS_BUSY[19][7] , 
        \ACCESS_BUSY[20][0] , \ACCESS_BUSY[20][1] , 
        \ACCESS_BUSY[20][2] , \ACCESS_BUSY[20][3] , 
        \ACCESS_BUSY[20][4] , \ACCESS_BUSY[20][5] , 
        \ACCESS_BUSY[20][6] , \ACCESS_BUSY[20][7] , 
        \ACCESS_BUSY[21][0] , \ACCESS_BUSY[21][1] , 
        \ACCESS_BUSY[21][2] , \ACCESS_BUSY[21][3] , 
        \ACCESS_BUSY[21][4] , \ACCESS_BUSY[21][5] , 
        \ACCESS_BUSY[21][6] , \ACCESS_BUSY[21][7] , 
        \ACCESS_BUSY[22][0] , \ACCESS_BUSY[22][1] , 
        \ACCESS_BUSY[22][2] , \ACCESS_BUSY[22][3] , 
        \ACCESS_BUSY[22][4] , \ACCESS_BUSY[22][5] , 
        \ACCESS_BUSY[22][6] , \ACCESS_BUSY[22][7] , 
        \ACCESS_BUSY[23][0] , \ACCESS_BUSY[23][1] , 
        \ACCESS_BUSY[23][2] , \ACCESS_BUSY[23][3] , 
        \ACCESS_BUSY[23][4] , \ACCESS_BUSY[23][5] , 
        \ACCESS_BUSY[23][6] , \ACCESS_BUSY[23][7] , 
        \ACCESS_BUSY[24][0] , \ACCESS_BUSY[24][1] , 
        \ACCESS_BUSY[24][2] , \ACCESS_BUSY[24][3] , 
        \ACCESS_BUSY[24][4] , \ACCESS_BUSY[24][5] , 
        \ACCESS_BUSY[24][6] , \ACCESS_BUSY[24][7] , 
        \ACCESS_BUSY[25][0] , \ACCESS_BUSY[25][1] , 
        \ACCESS_BUSY[25][2] , \ACCESS_BUSY[25][3] , 
        \ACCESS_BUSY[25][4] , \ACCESS_BUSY[25][5] , 
        \ACCESS_BUSY[25][6] , \ACCESS_BUSY[25][7] , 
        \ACCESS_BUSY[26][0] , \ACCESS_BUSY[26][1] , 
        \ACCESS_BUSY[26][2] , \ACCESS_BUSY[26][3] , 
        \ACCESS_BUSY[26][4] , \ACCESS_BUSY[26][5] , 
        \ACCESS_BUSY[26][6] , \ACCESS_BUSY[26][7] , 
        \ACCESS_BUSY[27][0] , \ACCESS_BUSY[27][1] , 
        \ACCESS_BUSY[27][2] , \ACCESS_BUSY[27][3] , 
        \ACCESS_BUSY[27][4] , \ACCESS_BUSY[27][5] , 
        \ACCESS_BUSY[27][6] , \ACCESS_BUSY[27][7] , 
        \ACCESS_BUSY[28][0] , \ACCESS_BUSY[28][1] , 
        \ACCESS_BUSY[28][2] , \ACCESS_BUSY[28][3] , 
        \ACCESS_BUSY[28][4] , \ACCESS_BUSY[28][5] , 
        \ACCESS_BUSY[28][6] , \ACCESS_BUSY[28][7] , 
        \ACCESS_BUSY[29][0] , \ACCESS_BUSY[29][1] , 
        \ACCESS_BUSY[29][2] , \ACCESS_BUSY[29][3] , 
        \ACCESS_BUSY[29][4] , \ACCESS_BUSY[29][5] , 
        \ACCESS_BUSY[29][6] , \ACCESS_BUSY[29][7] , 
        \ACCESS_BUSY[30][0] , \ACCESS_BUSY[30][1] , 
        \ACCESS_BUSY[30][2] , \ACCESS_BUSY[30][3] , 
        \ACCESS_BUSY[30][4] , \ACCESS_BUSY[30][5] , 
        \ACCESS_BUSY[30][6] , \ACCESS_BUSY[30][7] , 
        \ACCESS_BUSY[31][0] , \ACCESS_BUSY[31][1] , 
        \ACCESS_BUSY[31][2] , \ACCESS_BUSY[31][3] , 
        \ACCESS_BUSY[31][4] , \ACCESS_BUSY[31][5] , 
        \ACCESS_BUSY[31][6] , \ACCESS_BUSY[31][7] , 
        \ACCESS_BUSY[32][0] , \ACCESS_BUSY[32][1] , 
        \ACCESS_BUSY[32][2] , \ACCESS_BUSY[32][3] , 
        \ACCESS_BUSY[32][4] , \ACCESS_BUSY[32][5] , 
        \ACCESS_BUSY[32][6] , \ACCESS_BUSY[32][7] , 
        \ACCESS_BUSY[33][0] , \ACCESS_BUSY[33][1] , 
        \ACCESS_BUSY[33][2] , \ACCESS_BUSY[33][3] , 
        \ACCESS_BUSY[33][4] , \ACCESS_BUSY[33][5] , 
        \ACCESS_BUSY[33][6] , \ACCESS_BUSY[33][7] , 
        \ACCESS_BUSY[34][0] , \ACCESS_BUSY[34][1] , 
        \ACCESS_BUSY[34][2] , \ACCESS_BUSY[34][3] , 
        \ACCESS_BUSY[34][4] , \ACCESS_BUSY[34][5] , 
        \ACCESS_BUSY[34][6] , \ACCESS_BUSY[34][7] , 
        \ACCESS_BUSY[35][0] , \ACCESS_BUSY[35][1] , 
        \ACCESS_BUSY[35][2] , \ACCESS_BUSY[35][3] , 
        \ACCESS_BUSY[35][4] , \ACCESS_BUSY[35][5] , 
        \ACCESS_BUSY[35][6] , \ACCESS_BUSY[35][7] , 
        \ACCESS_BUSY[36][0] , \ACCESS_BUSY[36][1] , 
        \ACCESS_BUSY[36][2] , \ACCESS_BUSY[36][3] , 
        \ACCESS_BUSY[36][4] , \ACCESS_BUSY[36][5] , 
        \ACCESS_BUSY[36][6] , \ACCESS_BUSY[36][7] , 
        \ACCESS_BUSY[37][0] , \ACCESS_BUSY[37][1] , 
        \ACCESS_BUSY[37][2] , \ACCESS_BUSY[37][3] , 
        \ACCESS_BUSY[37][4] , \ACCESS_BUSY[37][5] , 
        \ACCESS_BUSY[37][6] , \ACCESS_BUSY[37][7] , 
        \ACCESS_BUSY[38][0] , \ACCESS_BUSY[38][1] , 
        \ACCESS_BUSY[38][2] , \ACCESS_BUSY[38][3] , 
        \ACCESS_BUSY[38][4] , \ACCESS_BUSY[38][5] , 
        \ACCESS_BUSY[38][6] , \ACCESS_BUSY[38][7] , 
        \ACCESS_BUSY[39][0] , \ACCESS_BUSY[39][1] , 
        \ACCESS_BUSY[39][2] , \ACCESS_BUSY[39][3] , 
        \ACCESS_BUSY[39][4] , \ACCESS_BUSY[39][5] , 
        \ACCESS_BUSY[39][6] , \ACCESS_BUSY[39][7] , 
        \ACCESS_BUSY[40][0] , \ACCESS_BUSY[40][1] , 
        \ACCESS_BUSY[40][2] , \ACCESS_BUSY[40][3] , 
        \ACCESS_BUSY[40][4] , \ACCESS_BUSY[40][5] , 
        \ACCESS_BUSY[40][6] , \ACCESS_BUSY[40][7] , 
        \ACCESS_BUSY[41][0] , \ACCESS_BUSY[41][1] , 
        \ACCESS_BUSY[41][2] , \ACCESS_BUSY[41][3] , 
        \ACCESS_BUSY[41][4] , \ACCESS_BUSY[41][5] , 
        \ACCESS_BUSY[41][6] , \ACCESS_BUSY[41][7] , 
        \ACCESS_BUSY[42][0] , \ACCESS_BUSY[42][1] , 
        \ACCESS_BUSY[42][2] , \ACCESS_BUSY[42][3] , 
        \ACCESS_BUSY[42][4] , \ACCESS_BUSY[42][5] , 
        \ACCESS_BUSY[42][6] , \ACCESS_BUSY[42][7] , 
        \ACCESS_BUSY[43][0] , \ACCESS_BUSY[43][1] , 
        \ACCESS_BUSY[43][2] , \ACCESS_BUSY[43][3] , 
        \ACCESS_BUSY[43][4] , \ACCESS_BUSY[43][5] , 
        \ACCESS_BUSY[43][6] , \ACCESS_BUSY[43][7] , 
        \ACCESS_BUSY[44][0] , \ACCESS_BUSY[44][1] , 
        \ACCESS_BUSY[44][2] , \ACCESS_BUSY[44][3] , 
        \ACCESS_BUSY[44][4] , \ACCESS_BUSY[44][5] , 
        \ACCESS_BUSY[44][6] , \ACCESS_BUSY[44][7] , 
        \ACCESS_BUSY[45][0] , \ACCESS_BUSY[45][1] , 
        \ACCESS_BUSY[45][2] , \ACCESS_BUSY[45][3] , 
        \ACCESS_BUSY[45][4] , \ACCESS_BUSY[45][5] , 
        \ACCESS_BUSY[45][6] , \ACCESS_BUSY[45][7] , 
        \ACCESS_BUSY[46][0] , \ACCESS_BUSY[46][1] , 
        \ACCESS_BUSY[46][2] , \ACCESS_BUSY[46][3] , 
        \ACCESS_BUSY[46][4] , \ACCESS_BUSY[46][5] , 
        \ACCESS_BUSY[46][6] , \ACCESS_BUSY[46][7] , 
        \ACCESS_BUSY[47][0] , \ACCESS_BUSY[47][1] , 
        \ACCESS_BUSY[47][2] , \ACCESS_BUSY[47][3] , 
        \ACCESS_BUSY[47][4] , \ACCESS_BUSY[47][5] , 
        \ACCESS_BUSY[47][6] , \ACCESS_BUSY[47][7] , 
        \ACCESS_BUSY[48][0] , \ACCESS_BUSY[48][1] , 
        \ACCESS_BUSY[48][2] , \ACCESS_BUSY[48][3] , 
        \ACCESS_BUSY[48][4] , \ACCESS_BUSY[48][5] , 
        \ACCESS_BUSY[48][6] , \ACCESS_BUSY[48][7] , 
        \ACCESS_BUSY[49][0] , \ACCESS_BUSY[49][1] , 
        \ACCESS_BUSY[49][2] , \ACCESS_BUSY[49][3] , 
        \ACCESS_BUSY[49][4] , \ACCESS_BUSY[49][5] , 
        \ACCESS_BUSY[49][6] , \ACCESS_BUSY[49][7] , 
        \ACCESS_BUSY[50][0] , \ACCESS_BUSY[50][1] , 
        \ACCESS_BUSY[50][2] , \ACCESS_BUSY[50][3] , 
        \ACCESS_BUSY[50][4] , \ACCESS_BUSY[50][5] , 
        \ACCESS_BUSY[50][6] , \ACCESS_BUSY[50][7] , 
        \ACCESS_BUSY[51][0] , \ACCESS_BUSY[51][1] , 
        \ACCESS_BUSY[51][2] , \ACCESS_BUSY[51][3] , 
        \ACCESS_BUSY[51][4] , \ACCESS_BUSY[51][5] , 
        \ACCESS_BUSY[51][6] , \ACCESS_BUSY[51][7] , 
        \ACCESS_BUSY[52][0] , \ACCESS_BUSY[52][1] , 
        \ACCESS_BUSY[52][2] , \ACCESS_BUSY[52][3] , 
        \ACCESS_BUSY[52][4] , \ACCESS_BUSY[52][5] , 
        \ACCESS_BUSY[52][6] , \ACCESS_BUSY[52][7] , 
        \ACCESS_BUSY[53][0] , \ACCESS_BUSY[53][1] , 
        \ACCESS_BUSY[53][2] , \ACCESS_BUSY[53][3] , 
        \ACCESS_BUSY[53][4] , \ACCESS_BUSY[53][5] , 
        \ACCESS_BUSY[53][6] , \ACCESS_BUSY[53][7] , 
        \ACCESS_BUSY[54][0] , \ACCESS_BUSY[54][1] , 
        \ACCESS_BUSY[54][2] , \ACCESS_BUSY[54][3] , 
        \ACCESS_BUSY[54][4] , \ACCESS_BUSY[54][5] , 
        \ACCESS_BUSY[54][6] , \ACCESS_BUSY[54][7] , 
        \ACCESS_BUSY[55][0] , \ACCESS_BUSY[55][1] , 
        \ACCESS_BUSY[55][2] , \ACCESS_BUSY[55][3] , 
        \ACCESS_BUSY[55][4] , \ACCESS_BUSY[55][5] , 
        \ACCESS_BUSY[55][6] , \ACCESS_BUSY[55][7] , 
        \ACCESS_BUSY[56][0] , \ACCESS_BUSY[56][1] , 
        \ACCESS_BUSY[56][2] , \ACCESS_BUSY[56][3] , 
        \ACCESS_BUSY[56][4] , \ACCESS_BUSY[56][5] , 
        \ACCESS_BUSY[56][6] , \ACCESS_BUSY[56][7] , 
        \ACCESS_BUSY[57][0] , \ACCESS_BUSY[57][1] , 
        \ACCESS_BUSY[57][2] , \ACCESS_BUSY[57][3] , 
        \ACCESS_BUSY[57][4] , \ACCESS_BUSY[57][5] , 
        \ACCESS_BUSY[57][6] , \ACCESS_BUSY[57][7] , 
        \ACCESS_BUSY[58][0] , \ACCESS_BUSY[58][1] , 
        \ACCESS_BUSY[58][2] , \ACCESS_BUSY[58][3] , 
        \ACCESS_BUSY[58][4] , \ACCESS_BUSY[58][5] , 
        \ACCESS_BUSY[58][6] , \ACCESS_BUSY[58][7] , 
        \ACCESS_BUSY[59][0] , \ACCESS_BUSY[59][1] , 
        \ACCESS_BUSY[59][2] , \ACCESS_BUSY[59][3] , 
        \ACCESS_BUSY[59][4] , \ACCESS_BUSY[59][5] , 
        \ACCESS_BUSY[59][6] , \ACCESS_BUSY[59][7] , 
        \ACCESS_BUSY[60][0] , \ACCESS_BUSY[60][1] , 
        \ACCESS_BUSY[60][2] , \ACCESS_BUSY[60][3] , 
        \ACCESS_BUSY[60][4] , \ACCESS_BUSY[60][5] , 
        \ACCESS_BUSY[60][6] , \ACCESS_BUSY[60][7] , 
        \ACCESS_BUSY[61][0] , \ACCESS_BUSY[61][1] , 
        \ACCESS_BUSY[61][2] , \ACCESS_BUSY[61][3] , 
        \ACCESS_BUSY[61][4] , \ACCESS_BUSY[61][5] , 
        \ACCESS_BUSY[61][6] , \ACCESS_BUSY[61][7] , 
        \ACCESS_BUSY[62][0] , \ACCESS_BUSY[62][1] , 
        \ACCESS_BUSY[62][2] , \ACCESS_BUSY[62][3] , 
        \ACCESS_BUSY[62][4] , \ACCESS_BUSY[62][5] , 
        \ACCESS_BUSY[62][6] , \ACCESS_BUSY[62][7] , 
        \ACCESS_BUSY[63][0] , \ACCESS_BUSY[63][1] , 
        \ACCESS_BUSY[63][2] , \ACCESS_BUSY[63][3] , 
        \ACCESS_BUSY[63][4] , \ACCESS_BUSY[63][5] , 
        \ACCESS_BUSY[63][6] , \ACCESS_BUSY[63][7] , 
        \ACCESS_BUSY[64][0] , \ACCESS_BUSY[64][1] , 
        \ACCESS_BUSY[64][2] , \ACCESS_BUSY[64][3] , 
        \ACCESS_BUSY[64][4] , \ACCESS_BUSY[64][5] , 
        \ACCESS_BUSY[64][6] , \ACCESS_BUSY[64][7] , 
        \ACCESS_BUSY[65][0] , \ACCESS_BUSY[65][1] , 
        \ACCESS_BUSY[65][2] , \ACCESS_BUSY[65][3] , 
        \ACCESS_BUSY[65][4] , \ACCESS_BUSY[65][5] , 
        \ACCESS_BUSY[65][6] , \ACCESS_BUSY[65][7] , 
        \ACCESS_BUSY[66][0] , \ACCESS_BUSY[66][1] , 
        \ACCESS_BUSY[66][2] , \ACCESS_BUSY[66][3] , 
        \ACCESS_BUSY[66][4] , \ACCESS_BUSY[66][5] , 
        \ACCESS_BUSY[66][6] , \ACCESS_BUSY[66][7] , 
        \ACCESS_BUSY[67][0] , \ACCESS_BUSY[67][1] , 
        \ACCESS_BUSY[67][2] , \ACCESS_BUSY[67][3] , 
        \ACCESS_BUSY[67][4] , \ACCESS_BUSY[67][5] , 
        \ACCESS_BUSY[67][6] , \ACCESS_BUSY[67][7] , 
        \ACCESS_BUSY[68][0] , \ACCESS_BUSY[68][1] , 
        \ACCESS_BUSY[68][2] , \ACCESS_BUSY[68][3] , 
        \ACCESS_BUSY[68][4] , \ACCESS_BUSY[68][5] , 
        \ACCESS_BUSY[68][6] , \ACCESS_BUSY[68][7] , 
        \ACCESS_BUSY[69][0] , \ACCESS_BUSY[69][1] , 
        \ACCESS_BUSY[69][2] , \ACCESS_BUSY[69][3] , 
        \ACCESS_BUSY[69][4] , \ACCESS_BUSY[69][5] , 
        \ACCESS_BUSY[69][6] , \ACCESS_BUSY[69][7] , 
        \ACCESS_BUSY[70][0] , \ACCESS_BUSY[70][1] , 
        \ACCESS_BUSY[70][2] , \ACCESS_BUSY[70][3] , 
        \ACCESS_BUSY[70][4] , \ACCESS_BUSY[70][5] , 
        \ACCESS_BUSY[70][6] , \ACCESS_BUSY[70][7] , 
        \ACCESS_BUSY[71][0] , \ACCESS_BUSY[71][1] , 
        \ACCESS_BUSY[71][2] , \ACCESS_BUSY[71][3] , 
        \ACCESS_BUSY[71][4] , \ACCESS_BUSY[71][5] , 
        \ACCESS_BUSY[71][6] , \ACCESS_BUSY[71][7] , 
        \ACCESS_BUSY[72][0] , \ACCESS_BUSY[72][1] , 
        \ACCESS_BUSY[72][2] , \ACCESS_BUSY[72][3] , 
        \ACCESS_BUSY[72][4] , \ACCESS_BUSY[72][5] , 
        \ACCESS_BUSY[72][6] , \ACCESS_BUSY[72][7] , 
        \ACCESS_BUSY[73][0] , \ACCESS_BUSY[73][1] , 
        \ACCESS_BUSY[73][2] , \ACCESS_BUSY[73][3] , 
        \ACCESS_BUSY[73][4] , \ACCESS_BUSY[73][5] , 
        \ACCESS_BUSY[73][6] , \ACCESS_BUSY[73][7] , 
        \ACCESS_BUSY[74][0] , \ACCESS_BUSY[74][1] , 
        \ACCESS_BUSY[74][2] , \ACCESS_BUSY[74][3] , 
        \ACCESS_BUSY[74][4] , \ACCESS_BUSY[74][5] , 
        \ACCESS_BUSY[74][6] , \ACCESS_BUSY[74][7] , 
        \ACCESS_BUSY[75][0] , \ACCESS_BUSY[75][1] , 
        \ACCESS_BUSY[75][2] , \ACCESS_BUSY[75][3] , 
        \ACCESS_BUSY[75][4] , \ACCESS_BUSY[75][5] , 
        \ACCESS_BUSY[75][6] , \ACCESS_BUSY[75][7] , 
        \ACCESS_BUSY[76][0] , \ACCESS_BUSY[76][1] , 
        \ACCESS_BUSY[76][2] , \ACCESS_BUSY[76][3] , 
        \ACCESS_BUSY[76][4] , \ACCESS_BUSY[76][5] , 
        \ACCESS_BUSY[76][6] , \ACCESS_BUSY[76][7] , 
        \ACCESS_BUSY[77][0] , \ACCESS_BUSY[77][1] , 
        \ACCESS_BUSY[77][2] , \ACCESS_BUSY[77][3] , 
        \ACCESS_BUSY[77][4] , \ACCESS_BUSY[77][5] , 
        \ACCESS_BUSY[77][6] , \ACCESS_BUSY[77][7] , 
        \ACCESS_BUSY[78][0] , \ACCESS_BUSY[78][1] , 
        \ACCESS_BUSY[78][2] , \ACCESS_BUSY[78][3] , 
        \ACCESS_BUSY[78][4] , \ACCESS_BUSY[78][5] , 
        \ACCESS_BUSY[78][6] , \ACCESS_BUSY[78][7] , 
        \ACCESS_BUSY[79][0] , \ACCESS_BUSY[79][1] , 
        \ACCESS_BUSY[79][2] , \ACCESS_BUSY[79][3] , 
        \ACCESS_BUSY[79][4] , \ACCESS_BUSY[79][5] , 
        \ACCESS_BUSY[79][6] , \ACCESS_BUSY[79][7] , 
        \ACCESS_BUSY[80][0] , \ACCESS_BUSY[80][1] , 
        \ACCESS_BUSY[80][2] , \ACCESS_BUSY[80][3] , 
        \ACCESS_BUSY[80][4] , \ACCESS_BUSY[80][5] , 
        \ACCESS_BUSY[80][6] , \ACCESS_BUSY[80][7] , 
        \ACCESS_BUSY[81][0] , \ACCESS_BUSY[81][1] , 
        \ACCESS_BUSY[81][2] , \ACCESS_BUSY[81][3] , 
        \ACCESS_BUSY[81][4] , \ACCESS_BUSY[81][5] , 
        \ACCESS_BUSY[81][6] , \ACCESS_BUSY[81][7] , 
        \ACCESS_BUSY[82][0] , \ACCESS_BUSY[82][1] , 
        \ACCESS_BUSY[82][2] , \ACCESS_BUSY[82][3] , 
        \ACCESS_BUSY[82][4] , \ACCESS_BUSY[82][5] , 
        \ACCESS_BUSY[82][6] , \ACCESS_BUSY[82][7] , 
        \ACCESS_BUSY[83][0] , \ACCESS_BUSY[83][1] , 
        \ACCESS_BUSY[83][2] , \ACCESS_BUSY[83][3] , 
        \ACCESS_BUSY[83][4] , \ACCESS_BUSY[83][5] , 
        \ACCESS_BUSY[83][6] , \ACCESS_BUSY[83][7] , 
        \ACCESS_BUSY[84][0] , \ACCESS_BUSY[84][1] , 
        \ACCESS_BUSY[84][2] , \ACCESS_BUSY[84][3] , 
        \ACCESS_BUSY[84][4] , \ACCESS_BUSY[84][5] , 
        \ACCESS_BUSY[84][6] , \ACCESS_BUSY[84][7] , 
        \ACCESS_BUSY[85][0] , \ACCESS_BUSY[85][1] , 
        \ACCESS_BUSY[85][2] , \ACCESS_BUSY[85][3] , 
        \ACCESS_BUSY[85][4] , \ACCESS_BUSY[85][5] , 
        \ACCESS_BUSY[85][6] , \ACCESS_BUSY[85][7] , 
        \ACCESS_BUSY[86][0] , \ACCESS_BUSY[86][1] , 
        \ACCESS_BUSY[86][2] , \ACCESS_BUSY[86][3] , 
        \ACCESS_BUSY[86][4] , \ACCESS_BUSY[86][5] , 
        \ACCESS_BUSY[86][6] , \ACCESS_BUSY[86][7] , 
        \ACCESS_BUSY[87][0] , \ACCESS_BUSY[87][1] , 
        \ACCESS_BUSY[87][2] , \ACCESS_BUSY[87][3] , 
        \ACCESS_BUSY[87][4] , \ACCESS_BUSY[87][5] , 
        \ACCESS_BUSY[87][6] , \ACCESS_BUSY[87][7] , 
        \ACCESS_BUSY[88][0] , \ACCESS_BUSY[88][1] , 
        \ACCESS_BUSY[88][2] , \ACCESS_BUSY[88][3] , 
        \ACCESS_BUSY[88][4] , \ACCESS_BUSY[88][5] , 
        \ACCESS_BUSY[88][6] , \ACCESS_BUSY[88][7] , 
        \ACCESS_BUSY[89][0] , \ACCESS_BUSY[89][1] , 
        \ACCESS_BUSY[89][2] , \ACCESS_BUSY[89][3] , 
        \ACCESS_BUSY[89][4] , \ACCESS_BUSY[89][5] , 
        \ACCESS_BUSY[89][6] , \ACCESS_BUSY[89][7] , 
        \ACCESS_BUSY[90][0] , \ACCESS_BUSY[90][1] , 
        \ACCESS_BUSY[90][2] , \ACCESS_BUSY[90][3] , 
        \ACCESS_BUSY[90][4] , \ACCESS_BUSY[90][5] , 
        \ACCESS_BUSY[90][6] , \ACCESS_BUSY[90][7] , 
        \ACCESS_BUSY[91][0] , \ACCESS_BUSY[91][1] , 
        \ACCESS_BUSY[91][2] , \ACCESS_BUSY[91][3] , 
        \ACCESS_BUSY[91][4] , \ACCESS_BUSY[91][5] , 
        \ACCESS_BUSY[91][6] , \ACCESS_BUSY[91][7] , 
        \ACCESS_BUSY[92][0] , \ACCESS_BUSY[92][1] , 
        \ACCESS_BUSY[92][2] , \ACCESS_BUSY[92][3] , 
        \ACCESS_BUSY[92][4] , \ACCESS_BUSY[92][5] , 
        \ACCESS_BUSY[92][6] , \ACCESS_BUSY[92][7] , 
        \ACCESS_BUSY[93][0] , \ACCESS_BUSY[93][1] , 
        \ACCESS_BUSY[93][2] , \ACCESS_BUSY[93][3] , 
        \ACCESS_BUSY[93][4] , \ACCESS_BUSY[93][5] , 
        \ACCESS_BUSY[93][6] , \ACCESS_BUSY[93][7] , 
        \ACCESS_BUSY[94][0] , \ACCESS_BUSY[94][1] , 
        \ACCESS_BUSY[94][2] , \ACCESS_BUSY[94][3] , 
        \ACCESS_BUSY[94][4] , \ACCESS_BUSY[94][5] , 
        \ACCESS_BUSY[94][6] , \ACCESS_BUSY[94][7] , 
        \ACCESS_BUSY[95][0] , \ACCESS_BUSY[95][1] , 
        \ACCESS_BUSY[95][2] , \ACCESS_BUSY[95][3] , 
        \ACCESS_BUSY[95][4] , \ACCESS_BUSY[95][5] , 
        \ACCESS_BUSY[95][6] , \ACCESS_BUSY[95][7] , 
        \ACCESS_BUSY[96][0] , \ACCESS_BUSY[96][1] , 
        \ACCESS_BUSY[96][2] , \ACCESS_BUSY[96][3] , 
        \ACCESS_BUSY[96][4] , \ACCESS_BUSY[96][5] , 
        \ACCESS_BUSY[96][6] , \ACCESS_BUSY[96][7] , 
        \ACCESS_BUSY[97][0] , \ACCESS_BUSY[97][1] , 
        \ACCESS_BUSY[97][2] , \ACCESS_BUSY[97][3] , 
        \ACCESS_BUSY[97][4] , \ACCESS_BUSY[97][5] , 
        \ACCESS_BUSY[97][6] , \ACCESS_BUSY[97][7] , 
        \ACCESS_BUSY[98][0] , \ACCESS_BUSY[98][1] , 
        \ACCESS_BUSY[98][2] , \ACCESS_BUSY[98][3] , 
        \ACCESS_BUSY[98][4] , \ACCESS_BUSY[98][5] , 
        \ACCESS_BUSY[98][6] , \ACCESS_BUSY[98][7] , 
        \ACCESS_BUSY[99][0] , \ACCESS_BUSY[99][1] , 
        \ACCESS_BUSY[99][2] , \ACCESS_BUSY[99][3] , 
        \ACCESS_BUSY[99][4] , \ACCESS_BUSY[99][5] , 
        \ACCESS_BUSY[99][6] , \ACCESS_BUSY[99][7] , 
        \ACCESS_BUSY[100][0] , \ACCESS_BUSY[100][1] , 
        \ACCESS_BUSY[100][2] , \ACCESS_BUSY[100][3] , 
        \ACCESS_BUSY[100][4] , \ACCESS_BUSY[100][5] , 
        \ACCESS_BUSY[100][6] , \ACCESS_BUSY[100][7] , 
        \ACCESS_BUSY[101][0] , \ACCESS_BUSY[101][1] , 
        \ACCESS_BUSY[101][2] , \ACCESS_BUSY[101][3] , 
        \ACCESS_BUSY[101][4] , \ACCESS_BUSY[101][5] , 
        \ACCESS_BUSY[101][6] , \ACCESS_BUSY[101][7] , 
        \ACCESS_BUSY[102][0] , \ACCESS_BUSY[102][1] , 
        \ACCESS_BUSY[102][2] , \ACCESS_BUSY[102][3] , 
        \ACCESS_BUSY[102][4] , \ACCESS_BUSY[102][5] , 
        \ACCESS_BUSY[102][6] , \ACCESS_BUSY[102][7] , 
        \ACCESS_BUSY[103][0] , \ACCESS_BUSY[103][1] , 
        \ACCESS_BUSY[103][2] , \ACCESS_BUSY[103][3] , 
        \ACCESS_BUSY[103][4] , \ACCESS_BUSY[103][5] , 
        \ACCESS_BUSY[103][6] , \ACCESS_BUSY[103][7] , 
        \ACCESS_BUSY[104][0] , \ACCESS_BUSY[104][1] , 
        \ACCESS_BUSY[104][2] , \ACCESS_BUSY[104][3] , 
        \ACCESS_BUSY[104][4] , \ACCESS_BUSY[104][5] , 
        \ACCESS_BUSY[104][6] , \ACCESS_BUSY[104][7] , 
        \ACCESS_BUSY[105][0] , \ACCESS_BUSY[105][1] , 
        \ACCESS_BUSY[105][2] , \ACCESS_BUSY[105][3] , 
        \ACCESS_BUSY[105][4] , \ACCESS_BUSY[105][5] , 
        \ACCESS_BUSY[105][6] , \ACCESS_BUSY[105][7] , 
        \ACCESS_BUSY[106][0] , \ACCESS_BUSY[106][1] , 
        \ACCESS_BUSY[106][2] , \ACCESS_BUSY[106][3] , 
        \ACCESS_BUSY[106][4] , \ACCESS_BUSY[106][5] , 
        \ACCESS_BUSY[106][6] , \ACCESS_BUSY[106][7] , 
        \ACCESS_BUSY[107][0] , \ACCESS_BUSY[107][1] , 
        \ACCESS_BUSY[107][2] , \ACCESS_BUSY[107][3] , 
        \ACCESS_BUSY[107][4] , \ACCESS_BUSY[107][5] , 
        \ACCESS_BUSY[107][6] , \ACCESS_BUSY[107][7] , 
        \ACCESS_BUSY[108][0] , \ACCESS_BUSY[108][1] , 
        \ACCESS_BUSY[108][2] , \ACCESS_BUSY[108][3] , 
        \ACCESS_BUSY[108][4] , \ACCESS_BUSY[108][5] , 
        \ACCESS_BUSY[108][6] , \ACCESS_BUSY[108][7] , 
        \ACCESS_BUSY[109][0] , \ACCESS_BUSY[109][1] , 
        \ACCESS_BUSY[109][2] , \ACCESS_BUSY[109][3] , 
        \ACCESS_BUSY[109][4] , \ACCESS_BUSY[109][5] , 
        \ACCESS_BUSY[109][6] , \ACCESS_BUSY[109][7] , 
        \ACCESS_BUSY[110][0] , \ACCESS_BUSY[110][1] , 
        \ACCESS_BUSY[110][2] , \ACCESS_BUSY[110][3] , 
        \ACCESS_BUSY[110][4] , \ACCESS_BUSY[110][5] , 
        \ACCESS_BUSY[110][6] , \ACCESS_BUSY[110][7] , 
        \ACCESS_BUSY[111][0] , \ACCESS_BUSY[111][1] , 
        \ACCESS_BUSY[111][2] , \ACCESS_BUSY[111][3] , 
        \ACCESS_BUSY[111][4] , \ACCESS_BUSY[111][5] , 
        \ACCESS_BUSY[111][6] , \ACCESS_BUSY[111][7] , 
        \ACCESS_BUSY[112][0] , \ACCESS_BUSY[112][1] , 
        \ACCESS_BUSY[112][2] , \ACCESS_BUSY[112][3] , 
        \ACCESS_BUSY[112][4] , \ACCESS_BUSY[112][5] , 
        \ACCESS_BUSY[112][6] , \ACCESS_BUSY[112][7] , 
        \ACCESS_BUSY[113][0] , \ACCESS_BUSY[113][1] , 
        \ACCESS_BUSY[113][2] , \ACCESS_BUSY[113][3] , 
        \ACCESS_BUSY[113][4] , \ACCESS_BUSY[113][5] , 
        \ACCESS_BUSY[113][6] , \ACCESS_BUSY[113][7] , 
        \ACCESS_BUSY[114][0] , \ACCESS_BUSY[114][1] , 
        \ACCESS_BUSY[114][2] , \ACCESS_BUSY[114][3] , 
        \ACCESS_BUSY[114][4] , \ACCESS_BUSY[114][5] , 
        \ACCESS_BUSY[114][6] , \ACCESS_BUSY[114][7] , 
        \ACCESS_BUSY[115][0] , \ACCESS_BUSY[115][1] , 
        \ACCESS_BUSY[115][2] , \ACCESS_BUSY[115][3] , 
        \ACCESS_BUSY[115][4] , \ACCESS_BUSY[115][5] , 
        \ACCESS_BUSY[115][6] , \ACCESS_BUSY[115][7] , 
        \ACCESS_BUSY[116][0] , \ACCESS_BUSY[116][1] , 
        \ACCESS_BUSY[116][2] , \ACCESS_BUSY[116][3] , 
        \ACCESS_BUSY[116][4] , \ACCESS_BUSY[116][5] , 
        \ACCESS_BUSY[116][6] , \ACCESS_BUSY[116][7] , 
        \ACCESS_BUSY[117][0] , \ACCESS_BUSY[117][1] , 
        \ACCESS_BUSY[117][2] , \ACCESS_BUSY[117][3] , 
        \ACCESS_BUSY[117][4] , \ACCESS_BUSY[117][5] , 
        \ACCESS_BUSY[117][6] , \ACCESS_BUSY[117][7] , 
        \ACCESS_BUSY[118][0] , \ACCESS_BUSY[118][1] , 
        \ACCESS_BUSY[118][2] , \ACCESS_BUSY[118][3] , 
        \ACCESS_BUSY[118][4] , \ACCESS_BUSY[118][5] , 
        \ACCESS_BUSY[118][6] , \ACCESS_BUSY[118][7] , OR4_1541_Y, 
        OR4_2173_Y, OR4_975_Y, OR4_989_Y, OR4_1215_Y, OR4_1794_Y, 
        OR4_184_Y, OR4_1161_Y, OR4_240_Y, OR4_1390_Y, OR4_2877_Y, 
        OR4_1392_Y, OR4_2190_Y, OR4_1254_Y, OR4_1441_Y, OR4_1269_Y, 
        OR4_2115_Y, OR4_263_Y, OR4_1331_Y, OR4_2033_Y, OR4_469_Y, 
        OR4_2034_Y, OR4_2876_Y, OR4_1888_Y, OR4_2091_Y, OR4_1895_Y, 
        OR4_2792_Y, OR4_944_Y, OR4_1964_Y, OR4_777_Y, OR4_2239_Y, 
        OR4_779_Y, OR4_1612_Y, OR4_644_Y, OR4_858_Y, OR4_659_Y, 
        OR4_1521_Y, OR4_2739_Y, OR2_23_Y, OR4_156_Y, OR4_394_Y, 
        OR4_1219_Y, OR4_2015_Y, OR4_2060_Y, OR4_1525_Y, OR4_2692_Y, 
        OR4_2870_Y, OR4_866_Y, OR4_2912_Y, OR4_542_Y, OR4_848_Y, 
        OR4_2434_Y, OR4_308_Y, OR4_3022_Y, OR4_1457_Y, OR4_2044_Y, 
        OR4_1857_Y, OR4_1795_Y, OR4_74_Y, OR4_760_Y, OR4_1090_Y, 
        OR4_2686_Y, OR4_550_Y, OR4_186_Y, OR4_1682_Y, OR4_2251_Y, 
        OR4_2083_Y, OR4_2036_Y, OR4_889_Y, OR4_1568_Y, OR4_1864_Y, 
        OR4_424_Y, OR4_1358_Y, OR4_1019_Y, OR4_2483_Y, OR4_42_Y, 
        OR4_2906_Y, OR2_73_Y, OR4_1137_Y, OR4_675_Y, OR4_2021_Y, 
        OR4_1010_Y, OR4_2819_Y, OR4_52_Y, OR4_2565_Y, OR4_616_Y, 
        OR4_1470_Y, OR4_791_Y, OR4_1480_Y, OR4_1775_Y, OR4_342_Y, 
        OR4_1282_Y, OR4_941_Y, OR4_2398_Y, OR4_3004_Y, OR4_2825_Y, 
        OR4_2775_Y, OR4_336_Y, OR4_1065_Y, OR4_1356_Y, OR4_2962_Y, 
        OR4_826_Y, OR4_468_Y, OR4_1963_Y, OR4_2544_Y, OR4_2350_Y, 
        OR4_2291_Y, OR4_1683_Y, OR4_2377_Y, OR4_2701_Y, OR4_1270_Y, 
        OR4_2150_Y, OR4_1809_Y, OR4_266_Y, OR4_869_Y, OR4_669_Y, 
        OR2_18_Y, OR4_2699_Y, OR4_429_Y, OR4_2400_Y, OR4_2195_Y, 
        OR4_2576_Y, OR4_360_Y, OR4_38_Y, OR4_1784_Y, OR4_2031_Y, 
        OR4_2019_Y, OR4_2659_Y, OR4_1831_Y, OR4_809_Y, OR4_1130_Y, 
        OR4_732_Y, OR4_1146_Y, OR4_1872_Y, OR4_2707_Y, OR4_1737_Y, 
        OR4_2832_Y, OR4_399_Y, OR4_2636_Y, OR4_1596_Y, OR4_1902_Y, 
        OR4_1533_Y, OR4_1925_Y, OR4_2678_Y, OR4_434_Y, OR4_2541_Y, 
        OR4_1731_Y, OR4_2367_Y, OR4_1565_Y, OR4_540_Y, OR4_852_Y, 
        OR4_474_Y, OR4_876_Y, OR4_1597_Y, OR4_2407_Y, OR2_35_Y, 
        OR4_2300_Y, OR4_901_Y, OR4_1830_Y, OR4_1501_Y, OR4_1993_Y, 
        OR4_2979_Y, OR4_2014_Y, OR4_521_Y, OR4_1108_Y, OR4_1632_Y, 
        OR4_2260_Y, OR4_1456_Y, OR4_428_Y, OR4_729_Y, OR4_369_Y, 
        OR4_750_Y, OR4_1495_Y, OR4_2304_Y, OR4_1387_Y, OR4_210_Y, 
        OR4_865_Y, OR4_47_Y, OR4_2048_Y, OR4_2343_Y, OR4_1982_Y, 
        OR4_2357_Y, OR4_73_Y, OR4_904_Y, OR4_3002_Y, OR4_1187_Y, 
        OR4_1792_Y, OR4_1011_Y, OR4_3010_Y, OR4_257_Y, OR4_2955_Y, 
        OR4_273_Y, OR4_1046_Y, OR4_1834_Y, OR2_27_Y, OR4_2690_Y, 
        OR4_3012_Y, OR4_800_Y, OR4_870_Y, OR4_2244_Y, OR4_2431_Y, 
        OR4_1362_Y, OR4_992_Y, OR4_1106_Y, OR4_2985_Y, OR4_2543_Y, 
        OR4_1198_Y, OR4_619_Y, OR4_1940_Y, OR4_1580_Y, OR4_2646_Y, 
        OR4_1314_Y, OR4_2749_Y, OR4_2193_Y, OR4_246_Y, OR4_2887_Y, 
        OR4_1494_Y, OR4_968_Y, OR4_2238_Y, OR4_1903_Y, OR4_2974_Y, 
        OR4_1614_Y, OR4_22_Y, OR4_2539_Y, OR4_1113_Y, OR4_670_Y, 
        OR4_2328_Y, OR4_1772_Y, OR4_61_Y, OR4_2768_Y, OR4_755_Y, 
        OR4_2459_Y, OR4_863_Y, OR2_9_Y, OR4_2689_Y, OR4_277_Y, 
        OR4_2078_Y, OR4_2093_Y, OR4_2308_Y, OR4_2950_Y, OR4_1337_Y, 
        OR4_2250_Y, OR4_1384_Y, OR4_2339_Y, OR4_21_Y, OR4_293_Y, 
        OR4_1906_Y, OR4_2847_Y, OR4_2463_Y, OR4_958_Y, OR4_1503_Y, 
        OR4_1340_Y, OR4_1283_Y, OR4_3009_Y, OR4_656_Y, OR4_973_Y, 
        OR4_2549_Y, OR4_425_Y, OR4_79_Y, OR4_1577_Y, OR4_2143_Y, 
        OR4_1967_Y, OR4_1911_Y, OR4_1742_Y, OR4_2438_Y, OR4_2765_Y, 
        OR4_1326_Y, OR4_2202_Y, OR4_1875_Y, OR4_323_Y, OR4_934_Y, 
        OR4_716_Y, OR2_21_Y, OR4_440_Y, OR4_2199_Y, OR4_1231_Y, 
        OR4_2378_Y, OR4_744_Y, OR4_219_Y, OR4_1553_Y, OR4_2480_Y, 
        OR4_2830_Y, OR4_271_Y, OR4_1751_Y, OR4_274_Y, OR4_1129_Y, 
        OR4_128_Y, OR4_330_Y, OR4_134_Y, OR4_1041_Y, OR4_2185_Y, 
        OR4_207_Y, OR4_2059_Y, OR4_502_Y, OR4_2063_Y, OR4_2919_Y, 
        OR4_1914_Y, OR4_2116_Y, OR4_1931_Y, OR4_2815_Y, OR4_972_Y, 
        OR4_1995_Y, OR4_1062_Y, OR4_2520_Y, OR4_1064_Y, OR4_1873_Y, 
        OR4_911_Y, OR4_1119_Y, OR4_928_Y, OR4_1769_Y, OR4_2982_Y, 
        OR2_30_Y, OR4_2335_Y, OR4_1165_Y, OR4_2771_Y, OR4_2120_Y, 
        OR4_768_Y, OR4_1919_Y, OR4_2263_Y, OR4_2744_Y, OR4_1044_Y, 
        OR4_1879_Y, OR4_1080_Y, OR4_6_Y, OR4_1637_Y, OR4_2648_Y, 
        OR4_278_Y, OR4_1952_Y, OR4_1346_Y, OR4_658_Y, OR4_2584_Y, 
        OR4_679_Y, OR4_2929_Y, OR4_1829_Y, OR4_450_Y, OR4_1439_Y, 
        OR4_2118_Y, OR4_741_Y, OR4_119_Y, OR4_2492_Y, OR4_1385_Y, 
        OR4_2262_Y, OR4_1454_Y, OR4_393_Y, OR4_2055_Y, OR4_20_Y, 
        OR4_688_Y, OR4_2340_Y, OR4_1714_Y, OR4_1077_Y, OR2_78_Y, 
        OR4_486_Y, OR4_75_Y, OR4_2814_Y, OR4_1718_Y, OR4_2081_Y, 
        OR4_2837_Y, OR4_2351_Y, OR4_1315_Y, OR4_2852_Y, OR4_298_Y, 
        OR4_1789_Y, OR4_301_Y, OR4_1167_Y, OR4_155_Y, OR4_375_Y, 
        OR4_170_Y, OR4_1074_Y, OR4_2220_Y, OR4_242_Y, OR4_2966_Y, 
        OR4_1395_Y, OR4_2968_Y, OR4_730_Y, OR4_2823_Y, OR4_3025_Y, 
        OR4_2839_Y, OR4_649_Y, OR4_1833_Y, OR4_2908_Y, OR4_2625_Y, 
        OR4_1084_Y, OR4_2631_Y, OR4_416_Y, OR4_2473_Y, OR4_2698_Y, 
        OR4_2486_Y, OR4_307_Y, OR4_1509_Y, OR2_65_Y, OR4_1761_Y, 
        OR4_1220_Y, OR4_935_Y, OR4_2401_Y, OR4_347_Y, OR4_2071_Y, 
        OR4_969_Y, OR4_1159_Y, OR4_738_Y, OR4_1116_Y, OR4_1719_Y, 
        OR4_950_Y, OR4_2953_Y, OR4_189_Y, OR4_2893_Y, OR4_203_Y, 
        OR4_979_Y, OR4_1764_Y, OR4_840_Y, OR4_529_Y, OR4_1185_Y, 
        OR4_338_Y, OR4_2353_Y, OR4_2679_Y, OR4_2282_Y, OR4_2695_Y, 
        OR4_385_Y, OR4_1225_Y, OR4_259_Y, OR4_235_Y, OR4_895_Y, 
        OR4_63_Y, OR4_2074_Y, OR4_2368_Y, OR4_2013_Y, OR4_2386_Y, 
        OR4_92_Y, OR4_943_Y, OR2_79_Y, OR4_439_Y, OR4_2754_Y, 
        OR4_2934_Y, OR4_1256_Y, OR4_593_Y, OR4_2980_Y, OR4_2484_Y, 
        OR4_2806_Y, OR4_175_Y, OR4_268_Y, OR4_1747_Y, OR4_270_Y, 
        OR4_1125_Y, OR4_126_Y, OR4_329_Y, OR4_132_Y, OR4_1039_Y, 
        OR4_2183_Y, OR4_201_Y, OR4_2569_Y, OR4_1031_Y, OR4_2574_Y, 
        OR4_352_Y, OR4_2410_Y, OR4_2632_Y, OR4_2422_Y, OR4_256_Y, 
        OR4_1446_Y, OR4_2499_Y, OR4_2761_Y, OR4_1203_Y, OR4_2763_Y, 
        OR4_539_Y, OR4_2610_Y, OR4_2828_Y, OR4_2618_Y, OR4_433_Y, 
        OR4_1625_Y, OR2_68_Y, OR4_2466_Y, OR4_605_Y, OR4_2333_Y, 
        OR4_1201_Y, OR4_2039_Y, OR4_1273_Y, OR4_1038_Y, OR4_522_Y, 
        OR4_497_Y, OR4_1798_Y, OR4_2430_Y, OR4_1617_Y, OR4_598_Y, 
        OR4_917_Y, OR4_535_Y, OR4_947_Y, OR4_1647_Y, OR4_2472_Y, 
        OR4_1536_Y, OR4_2992_Y, OR4_569_Y, OR4_2816_Y, OR4_1760_Y, 
        OR4_2073_Y, OR4_1692_Y, OR4_2090_Y, OR4_2859_Y, OR4_611_Y, 
        OR4_2732_Y, OR4_1668_Y, OR4_2297_Y, OR4_1487_Y, OR4_472_Y, 
        OR4_766_Y, OR4_401_Y, OR4_782_Y, OR4_1531_Y, OR4_2338_Y, 
        OR2_33_Y, OR4_1469_Y, OR4_501_Y, OR4_348_Y, OR4_125_Y, OR4_9_Y, 
        OR4_1589_Y, OR4_2809_Y, OR4_2506_Y, OR4_1640_Y, OR4_808_Y, 
        OR4_1440_Y, OR4_631_Y, OR4_2650_Y, OR4_2964_Y, OR4_2587_Y, 
        OR4_2977_Y, OR4_668_Y, OR4_1473_Y, OR4_544_Y, OR4_2892_Y, 
        OR4_466_Y, OR4_2704_Y, OR4_1646_Y, OR4_1962_Y, OR4_1588_Y, 
        OR4_1976_Y, OR4_2748_Y, OR4_506_Y, OR4_2612_Y, OR4_2751_Y, 
        OR4_309_Y, OR4_2546_Y, OR4_1517_Y, OR4_1815_Y, OR4_1447_Y, 
        OR4_1835_Y, OR4_2598_Y, OR4_356_Y, OR2_61_Y, OR4_2265_Y, 
        OR4_1235_Y, OR4_2700_Y, OR4_2169_Y, OR4_844_Y, OR4_1978_Y, 
        OR4_2330_Y, OR4_2666_Y, OR4_1101_Y, OR4_1808_Y, OR4_1021_Y, 
        OR4_2983_Y, OR4_1583_Y, OR4_2590_Y, OR4_213_Y, OR4_1889_Y, 
        OR4_1277_Y, OR4_592_Y, OR4_2508_Y, OR4_731_Y, OR4_2978_Y, 
        OR4_1899_Y, OR4_520_Y, OR4_1499_Y, OR4_2168_Y, OR4_815_Y, 
        OR4_179_Y, OR4_2554_Y, OR4_1434_Y, OR4_2191_Y, OR4_1406_Y, 
        OR4_325_Y, OR4_1990_Y, OR4_2994_Y, OR4_623_Y, OR4_2270_Y, 
        OR4_1656_Y, OR4_1017_Y, OR2_75_Y, OR4_2628_Y, OR4_2491_Y, 
        OR4_1648_Y, OR4_2266_Y, OR4_2296_Y, OR4_1333_Y, OR4_2249_Y, 
        OR4_437_Y, OR4_733_Y, OR4_1955_Y, OR4_2602_Y, OR4_1763_Y, 
        OR4_736_Y, OR4_1072_Y, OR4_681_Y, OR4_1091_Y, OR4_1804_Y, 
        OR4_2633_Y, OR4_1676_Y, OR4_1818_Y, OR4_2453_Y, OR4_1631_Y, 
        OR4_618_Y, OR4_951_Y, OR4_555_Y, OR4_963_Y, OR4_1672_Y, 
        OR4_2496_Y, OR4_1555_Y, OR4_1018_Y, OR4_1620_Y, OR4_814_Y, 
        OR4_2848_Y, OR4_84_Y, OR4_2787_Y, OR4_100_Y, OR4_862_Y, 
        OR4_1655_Y, OR2_24_Y, OR4_1956_Y, OR4_2665_Y, OR4_2404_Y, 
        OR4_1687_Y, OR4_1776_Y, OR4_603_Y, OR4_131_Y, OR4_2206_Y, 
        OR4_2921_Y, OR4_2225_Y, OR4_1814_Y, OR4_455_Y, OR4_2957_Y, 
        OR4_1239_Y, OR4_878_Y, OR4_1910_Y, OR4_578_Y, OR4_2004_Y, 
        OR4_1488_Y, OR4_2971_Y, OR4_2522_Y, OR4_1179_Y, OR4_597_Y, 
        OR4_1918_Y, OR4_1560_Y, OR4_2622_Y, OR4_1293_Y, OR4_2725_Y, 
        OR4_2174_Y, OR4_2733_Y, OR4_2264_Y, OR4_946_Y, OR4_351_Y, 
        OR4_1670_Y, OR4_1338_Y, OR4_2363_Y, OR4_1063_Y, OR4_2456_Y, 
        OR2_48_Y, OR4_1380_Y, OR4_16_Y, OR4_2946_Y, OR4_1458_Y, 
        OR4_715_Y, OR4_1713_Y, OR4_1216_Y, OR4_1559_Y, OR4_1601_Y, 
        OR4_916_Y, OR4_80_Y, OR4_2058_Y, OR4_678_Y, OR4_1650_Y, 
        OR4_2332_Y, OR4_995_Y, OR4_339_Y, OR4_2741_Y, OR4_1593_Y, 
        OR4_2581_Y, OR4_1743_Y, OR4_693_Y, OR4_2336_Y, OR4_287_Y, 
        OR4_1002_Y, OR4_2652_Y, OR4_2024_Y, OR4_1363_Y, OR4_224_Y, 
        OR4_2450_Y, OR4_1627_Y, OR4_571_Y, OR4_2205_Y, OR4_166_Y, 
        OR4_880_Y, OR4_2533_Y, OR4_1905_Y, OR4_1252_Y, OR2_2_Y, 
        OR4_1575_Y, OR4_297_Y, OR4_2318_Y, OR4_480_Y, OR4_1880_Y, 
        OR4_1365_Y, OR4_2697_Y, OR4_573_Y, OR4_909_Y, OR4_1266_Y, 
        OR4_1944_Y, OR4_2215_Y, OR4_804_Y, OR4_1706_Y, OR4_1379_Y, 
        OR4_2886_Y, OR4_403_Y, OR4_211_Y, OR4_150_Y, OR4_3039_Y, 
        OR4_685_Y, OR4_1005_Y, OR4_2600_Y, OR4_463_Y, OR4_104_Y, 
        OR4_1599_Y, OR4_2166_Y, OR4_1999_Y, OR4_1947_Y, OR4_2010_Y, 
        OR4_2724_Y, OR4_3014_Y, OR4_1567_Y, OR4_2476_Y, OR4_2125_Y, 
        OR4_589_Y, OR4_1190_Y, OR4_1004_Y, OR2_28_Y, OR4_1603_Y, 
        OR4_1226_Y, OR4_891_Y, OR4_2879_Y, OR4_153_Y, OR4_920_Y, 
        OR4_443_Y, OR4_2418_Y, OR4_940_Y, OR4_1297_Y, OR4_1975_Y, 
        OR4_2256_Y, OR4_854_Y, OR4_1754_Y, OR4_1410_Y, OR4_2931_Y, 
        OR4_438_Y, OR4_247_Y, OR4_192_Y, OR4_892_Y, OR4_1573_Y, 
        OR4_1869_Y, OR4_426_Y, OR4_1364_Y, OR4_1025_Y, OR4_2493_Y, 
        OR4_45_Y, OR4_2913_Y, OR4_2860_Y, OR4_554_Y, OR4_1263_Y, 
        OR4_1539_Y, OR4_103_Y, OR4_1049_Y, OR4_676_Y, OR4_2151_Y, 
        OR4_2772_Y, OR4_2562_Y, OR2_64_Y, OR4_1825_Y, OR4_2064_Y, 
        OR4_2873_Y, OR4_636_Y, OR4_680_Y, OR4_135_Y, OR4_1312_Y, 
        OR4_1468_Y, OR4_2510_Y, OR4_1184_Y, OR4_1791_Y, OR4_1009_Y, 
        OR4_3008_Y, OR4_254_Y, OR4_2951_Y, OR4_269_Y, OR4_1043_Y, 
        OR4_1832_Y, OR4_913_Y, OR4_1399_Y, OR4_2029_Y, OR4_1234_Y, 
        OR4_169_Y, OR4_491_Y, OR4_112_Y, OR4_508_Y, OR4_1267_Y, 
        OR4_2067_Y, OR4_1144_Y, OR4_2170_Y, OR4_2843_Y, OR4_2008_Y, 
        OR4_1007_Y, OR4_1298_Y, OR4_942_Y, OR4_1316_Y, OR4_2043_Y, 
        OR4_2878_Y, OR2_46_Y, OR4_2804_Y, OR4_2316_Y, OR4_642_Y, 
        OR4_2655_Y, OR4_1421_Y, OR4_1695_Y, OR4_1202_Y, OR4_2253_Y, 
        OR4_91_Y, OR4_2105_Y, OR4_2766_Y, OR4_1933_Y, OR4_921_Y, 
        OR4_1230_Y, OR4_846_Y, OR4_1244_Y, OR4_1968_Y, OR4_2810_Y, 
        OR4_1840_Y, OR4_1651_Y, OR4_2283_Y, OR4_1475_Y, OR4_453_Y, 
        OR4_752_Y, OR4_389_Y, OR4_770_Y, OR4_1519_Y, OR4_2321_Y, 
        OR4_1404_Y, OR4_3026_Y, OR4_606_Y, OR4_2855_Y, OR4_1796_Y, 
        OR4_2101_Y, OR4_1724_Y, OR4_2119_Y, OR4_2894_Y, OR4_647_Y, 
        OR2_70_Y, OR4_1571_Y, OR4_824_Y, OR4_1024_Y, OR4_2355_Y, 
        OR4_1701_Y, OR4_1076_Y, OR4_575_Y, OR4_882_Y, OR4_1330_Y, 
        OR4_1260_Y, OR4_1942_Y, OR4_2209_Y, OR4_801_Y, OR4_1704_Y, 
        OR4_1376_Y, OR4_2884_Y, OR4_400_Y, OR4_208_Y, OR4_148_Y, 
        OR4_495_Y, OR4_1206_Y, OR4_1478_Y, OR4_53_Y, OR4_986_Y, 
        OR4_615_Y, OR4_2104_Y, OR4_2709_Y, OR4_2504_Y, OR4_2439_Y, 
        OR4_674_Y, OR4_1377_Y, OR4_1653_Y, OR4_223_Y, OR4_1160_Y, 
        OR4_788_Y, OR4_2273_Y, OR4_2895_Y, OR4_2696_Y, OR2_66_Y, 
        OR4_1635_Y, OR4_29_Y, OR4_1087_Y, OR4_902_Y, OR4_2585_Y, 
        OR4_1355_Y, OR4_990_Y, OR4_2406_Y, OR4_1666_Y, OR4_1950_Y, 
        OR4_1515_Y, OR4_140_Y, OR4_2640_Y, OR4_937_Y, OR4_558_Y, 
        OR4_1604_Y, OR4_267_Y, OR4_1688_Y, OR4_1210_Y, OR4_294_Y, 
        OR4_2941_Y, OR4_1550_Y, OR4_1020_Y, OR4_2302_Y, OR4_1959_Y, 
        OR4_3028_Y, OR4_1669_Y, OR4_60_Y, OR4_2607_Y, OR4_1370_Y, 
        OR4_959_Y, OR4_2615_Y, OR4_2042_Y, OR4_312_Y, OR4_3023_Y, 
        OR4_1048_Y, OR4_2753_Y, OR4_1132_Y, OR2_17_Y, OR4_30_Y, 
        OR4_2326_Y, OR4_1755_Y, OR4_2164_Y, OR4_2113_Y, OR4_368_Y, 
        OR4_83_Y, OR4_707_Y, OR4_2163_Y, OR4_2911_Y, OR4_1345_Y, 
        OR4_2914_Y, OR4_682_Y, OR4_2762_Y, OR4_2969_Y, OR4_2783_Y, 
        OR4_587_Y, OR4_1767_Y, OR4_2844_Y, OR4_2155_Y, OR4_613_Y, 
        OR4_2156_Y, OR4_3021_Y, OR4_2035_Y, OR4_2208_Y, OR4_2041_Y, 
        OR4_2935_Y, OR4_1086_Y, OR4_2103_Y, OR4_1584_Y, OR4_40_Y, 
        OR4_1585_Y, OR4_2415_Y, OR4_1442_Y, OR4_1638_Y, OR4_1452_Y, 
        OR4_2311_Y, OR4_483_Y, OR2_38_Y, CFG3_11_Y, CFG3_8_Y, 
        CFG3_22_Y, CFG3_20_Y, CFG3_12_Y, CFG3_6_Y, CFG3_19_Y, CFG3_2_Y, 
        CFG3_16_Y, CFG3_15_Y, CFG3_21_Y, CFG3_9_Y, OR4_2820_Y, 
        OR4_255_Y, OR4_2495_Y, OR4_296_Y, OR4_1246_Y, OR4_2158_Y, 
        OR4_1342_Y, OR4_1649_Y, OR4_212_Y, OR4_2641_Y, OR4_1093_Y, 
        OR4_2642_Y, OR4_420_Y, OR4_2481_Y, OR4_2714_Y, OR4_2502_Y, 
        OR4_321_Y, OR4_1520_Y, OR4_2579_Y, OR4_87_Y, OR4_1576_Y, 
        OR4_88_Y, OR4_956_Y, OR4_3000_Y, OR4_143_Y, OR4_3016_Y, 
        OR4_835_Y, OR4_2026_Y, OR4_41_Y, OR4_2312_Y, OR4_761_Y, 
        OR4_2313_Y, OR4_118_Y, OR4_2165_Y, OR4_2380_Y, OR4_2175_Y, 
        OR4_37_Y, OR4_1241_Y, OR2_52_Y, OR4_945_Y, OR4_974_Y, 
        OR4_1214_Y, OR4_2807_Y, OR4_2525_Y, OR4_382_Y, OR4_1152_Y, 
        OR4_2677_Y, OR4_454_Y, OR4_1236_Y, OR4_776_Y, OR4_2452_Y, 
        OR4_1900_Y, OR4_165_Y, OR4_2883_Y, OR4_893_Y, OR4_2597_Y, 
        OR4_987_Y, OR4_460_Y, OR4_1265_Y, OR4_823_Y, OR4_2489_Y, 
        OR4_1936_Y, OR4_205_Y, OR4_2925_Y, OR4_933_Y, OR4_2621_Y, 
        OR4_1030_Y, OR4_498_Y, OR4_1481_Y, OR4_1082_Y, OR4_2759_Y, 
        OR4_2157_Y, OR4_456_Y, OR4_93_Y, OR4_1177_Y, OR4_2875_Y, 
        OR4_1258_Y, OR2_25_Y, OR4_1785_Y, OR4_1343_Y, OR4_2416_Y, 
        OR4_2374_Y, OR4_1036_Y, OR4_1974_Y, OR4_1276_Y, OR4_988_Y, 
        OR4_2097_Y, OR4_2089_Y, OR4_1644_Y, OR4_289_Y, OR4_2802_Y, 
        OR4_1078_Y, OR4_703_Y, OR4_1741_Y, OR4_418_Y, OR4_1836_Y, 
        OR4_1352_Y, OR4_1613_Y, OR4_1208_Y, OR4_2891_Y, OR4_2292_Y, 
        OR4_590_Y, OR4_226_Y, OR4_1299_Y, OR4_2999_Y, OR4_1383_Y, 
        OR4_883_Y, OR4_2747_Y, OR4_2278_Y, OR4_957_Y, OR4_364_Y, 
        OR4_1679_Y, OR4_1351_Y, OR4_2373_Y, OR4_1073_Y, OR4_2469_Y, 
        OR2_49_Y, OR4_1407_Y, OR4_1098_Y, OR4_967_Y, OR4_57_Y, 
        OR4_576_Y, OR4_1514_Y, OR4_317_Y, OR4_2419_Y, OR4_2216_Y, 
        OR4_1247_Y, OR4_2734_Y, OR4_1250_Y, OR4_2068_Y, OR4_1104_Y, 
        OR4_1306_Y, OR4_1117_Y, OR4_1970_Y, OR4_117_Y, OR4_1191_Y, 
        OR4_936_Y, OR4_2382_Y, OR4_938_Y, OR4_1735_Y, OR4_764_Y, 
        OR4_1001_Y, OR4_775_Y, OR4_1636_Y, OR4_2866_Y, OR4_864_Y, 
        OR4_765_Y, OR4_2227_Y, OR4_767_Y, OR4_1600_Y, OR4_632_Y, 
        OR4_841_Y, OR4_643_Y, OR4_1505_Y, OR4_2721_Y, OR2_22_Y, 
        OR4_1309_Y, OR4_1946_Y, OR4_704_Y, OR4_711_Y, OR4_970_Y, 
        OR4_1543_Y, OR4_2995_Y, OR4_907_Y, OR4_11_Y, OR4_628_Y, 
        OR4_1275_Y, OR4_442_Y, OR4_2454_Y, OR4_2790_Y, OR4_2384_Y, 
        OR4_2805_Y, OR4_489_Y, OR4_1313_Y, OR4_361_Y, OR4_1287_Y, 
        OR4_1907_Y, OR4_1110_Y, OR4_65_Y, OR4_366_Y, OR4_15_Y, 
        OR4_386_Y, OR4_1147_Y, OR4_1951_Y, OR4_1034_Y, OR4_39_Y, 
        OR4_667_Y, OR4_2917_Y, OR4_1862_Y, OR4_2149_Y, OR4_1790_Y, 
        OR4_2162_Y, OR4_2944_Y, OR4_705_Y, OR2_72_Y, OR4_2713_Y, 
        OR4_319_Y, OR4_349_Y, OR4_754_Y, OR4_313_Y, OR4_1408_Y, 
        OR4_3006_Y, OR4_372_Y, OR4_1781_Y, OR4_3001_Y, OR4_2563_Y, 
        OR4_1218_Y, OR4_638_Y, OR4_1958_Y, OR4_1595_Y, OR4_2663_Y, 
        OR4_1332_Y, OR4_2764_Y, OR4_2211_Y, OR4_625_Y, OR4_188_Y, 
        OR4_1871_Y, OR4_1327_Y, OR4_2639_Y, OR4_2255_Y, OR4_280_Y, 
        OR4_1994_Y, OR4_376_Y, OR4_2936_Y, OR4_655_Y, OR4_216_Y, 
        OR4_1898_Y, OR4_1353_Y, OR4_2670_Y, OR4_2290_Y, OR4_299_Y, 
        OR4_2020_Y, OR4_402_Y, OR2_77_Y, OR4_1158_Y, OR4_421_Y, 
        OR4_2909_Y, OR4_265_Y, OR4_197_Y, OR4_1491_Y, OR4_1237_Y, 
        OR4_1828_Y, OR4_264_Y, OR4_821_Y, OR4_1507_Y, OR4_1800_Y, 
        OR4_371_Y, OR4_1302_Y, OR4_961_Y, OR4_2424_Y, OR4_3030_Y, 
        OR4_2849_Y, OR4_2801_Y, OR4_97_Y, OR4_794_Y, OR4_1111_Y, 
        OR4_2718_Y, OR4_572_Y, OR4_217_Y, OR4_1705_Y, OR4_2289_Y, 
        OR4_2106_Y, OR4_2062_Y, OR4_2557_Y, OR4_206_Y, OR4_514_Y, 
        OR4_2109_Y, OR4_8_Y, OR4_2693_Y, OR4_1154_Y, OR4_1703_Y, 
        OR4_1528_Y, OR2_34_Y, OR4_925_Y, OR4_121_Y, OR4_1690_Y, 
        OR4_2824_Y, OR4_2811_Y, OR4_1986_Y, OR4_1422_Y, OR4_896_Y, 
        OR4_1_Y, OR4_430_Y, OR4_2673_Y, OR4_1587_Y, OR4_202_Y, 
        OR4_1221_Y, OR4_1887_Y, OR4_513_Y, OR4_2947_Y, OR4_2232_Y, 
        OR4_1149_Y, OR4_2720_Y, OR4_1884_Y, OR4_820_Y, OR4_2468_Y, 
        OR4_419_Y, OR4_1122_Y, OR4_2799_Y, OR4_2137_Y, OR4_1466_Y, 
        OR4_353_Y, OR4_1251_Y, OR4_415_Y, OR4_2375_Y, OR4_1033_Y, 
        OR4_1996_Y, OR4_2691_Y, OR4_1318_Y, OR4_684_Y, OR4_23_Y, 
        OR2_47_Y, OR4_2293_Y, OR4_236_Y, OR4_350_Y, OR4_231_Y, 
        OR4_2735_Y, OR4_620_Y, OR4_1115_Y, OR4_1842_Y, OR4_723_Y, 
        OR4_2132_Y, OR4_581_Y, OR4_2133_Y, OR4_2987_Y, OR4_1998_Y, 
        OR4_2180_Y, OR4_2011_Y, OR4_2903_Y, OR4_1052_Y, OR4_2076_Y, 
        OR4_76_Y, OR4_1551_Y, OR4_78_Y, OR4_930_Y, OR4_2986_Y, 
        OR4_129_Y, OR4_2996_Y, OR4_818_Y, OR4_2007_Y, OR4_28_Y, 
        OR4_173_Y, OR4_1658_Y, OR4_176_Y, OR4_1045_Y, OR4_50_Y, 
        OR4_241_Y, OR4_59_Y, OR4_955_Y, OR4_2111_Y, OR2_3_Y, 
        OR4_1782_Y, OR4_396_Y, OR4_580_Y, OR4_1817_Y, OR4_423_Y, 
        OR4_727_Y, OR4_570_Y, OR4_1109_Y, OR4_2395_Y, OR4_1615_Y, 
        OR4_62_Y, OR4_1616_Y, OR4_2448_Y, OR4_1471_Y, OR4_1673_Y, 
        OR4_1485_Y, OR4_2354_Y, OR4_515_Y, OR4_1558_Y, OR4_227_Y, 
        OR4_1699_Y, OR4_229_Y, OR4_1092_Y, OR4_85_Y, OR4_286_Y, 
        OR4_95_Y, OR4_994_Y, OR4_2147_Y, OR4_152_Y, OR4_412_Y, 
        OR4_1891_Y, OR4_414_Y, OR4_1264_Y, OR4_262_Y, OR4_476_Y, 
        OR4_275_Y, OR4_1169_Y, OR4_2327_Y, OR2_11_Y, OR4_903_Y, 
        OR4_1397_Y, OR4_585_Y, OR4_1433_Y, OR4_2349_Y, OR4_258_Y, 
        OR4_2443_Y, OR4_2813_Y, OR4_1360_Y, OR4_562_Y, OR4_1271_Y, 
        OR4_1549_Y, OR4_115_Y, OR4_1058_Y, OR4_687_Y, OR4_2160_Y, 
        OR4_2788_Y, OR4_2580_Y, OR4_2519_Y, OR4_1085_Y, OR4_1750_Y, 
        OR4_2054_Y, OR4_621_Y, OR4_1534_Y, OR4_1205_Y, OR4_2694_Y, 
        OR4_215_Y, OR4_44_Y, OR4_3033_Y, OR4_253_Y, OR4_976_Y, 
        OR4_1268_Y, OR4_2871_Y, OR4_722_Y, OR4_378_Y, OR4_1877_Y, 
        OR4_2447_Y, OR4_2247_Y, OR2_51_Y, OR4_2527_Y, OR4_2187_Y, 
        OR4_2069_Y, OR4_1200_Y, OR4_1693_Y, OR4_2654_Y, OR4_1448_Y, 
        OR4_519_Y, OR4_315_Y, OR4_2178_Y, OR4_2922_Y, OR4_139_Y, 
        OR4_1753_Y, OR4_2688_Y, OR4_2305_Y, OR4_773_Y, OR4_1371_Y, 
        OR4_1194_Y, OR4_1135_Y, OR4_1885_Y, OR4_2591_Y, OR4_2900_Y, 
        OR4_1435_Y, OR4_2348_Y, OR4_2006_Y, OR4_462_Y, OR4_1066_Y, 
        OR4_868_Y, OR4_797_Y, OR4_1729_Y, OR4_2426_Y, OR4_2756_Y, 
        OR4_1311_Y, OR4_2189_Y, OR4_1861_Y, OR4_304_Y, OR4_915_Y, 
        OR4_710_Y, OR2_19_Y, OR4_180_Y, OR4_1971_Y, OR4_977_Y, 
        OR4_2130_Y, OR4_504_Y, OR4_3027_Y, OR4_1317_Y, OR4_2210_Y, 
        OR4_2550_Y, OR4_2572_Y, OR4_144_Y, OR4_2372_Y, OR4_1368_Y, 
        OR4_1643_Y, OR4_1304_Y, OR4_1667_Y, OR4_2411_Y, OR4_190_Y, 
        OR4_2284_Y, OR4_1319_Y, OR4_1939_Y, OR4_1143_Y, OR4_89_Y, 
        OR4_397_Y, OR4_43_Y, OR4_417_Y, OR4_1182_Y, OR4_1972_Y, 
        OR4_1060_Y, OR4_279_Y, OR4_948_Y, OR4_99_Y, OR4_2112_Y, 
        OR4_2413_Y, OR4_2052_Y, OR4_2428_Y, OR4_130_Y, OR4_980_Y, 
        OR2_0_Y, OR4_225_Y, OR4_2882_Y, OR4_2537_Y, OR4_1474_Y, 
        OR4_1822_Y, OR4_2568_Y, OR4_2102_Y, OR4_1070_Y, OR4_2586_Y, 
        OR4_2611_Y, OR4_187_Y, OR4_2412_Y, OR4_1400_Y, OR4_1684_Y, 
        OR4_1348_Y, OR4_1700_Y, OR4_2449_Y, OR4_230_Y, OR4_2319_Y, 
        OR4_2172_Y, OR4_2851_Y, OR4_2017_Y, OR4_1012_Y, OR4_1303_Y, 
        OR4_952_Y, OR4_1323_Y, OR4_2049_Y, OR4_2890_Y, OR4_1930_Y, 
        OR4_1868_Y, OR4_2503_Y, OR4_1678_Y, OR4_665_Y, OR4_984_Y, 
        OR4_596_Y, OR4_1006_Y, OR4_1709_Y, OR4_2538_Y, OR2_39_Y, 
        OR4_1096_Y, OR4_792_Y, OR4_2942_Y, OR4_493_Y, OR4_1758_Y, 
        OR4_2131_Y, OR4_1732_Y, OR4_2784_Y, OR4_49_Y, OR4_929_Y, 
        OR4_2376_Y, OR4_932_Y, OR4_1730_Y, OR4_758_Y, OR4_998_Y, 
        OR4_772_Y, OR4_1634_Y, OR4_2864_Y, OR4_856_Y, OR4_626_Y, 
        OR4_2099_Y, OR4_630_Y, OR4_1453_Y, OR4_488_Y, OR4_695_Y, 
        OR4_500_Y, OR4_1375_Y, OR4_2553_Y, OR4_563_Y, OR4_2780_Y, 
        OR4_1209_Y, OR4_2782_Y, OR4_551_Y, OR4_2617_Y, OR4_2838_Y, 
        OR4_2629_Y, OR4_449_Y, OR4_1630_Y, OR2_69_Y, OR4_641_Y, 
        OR4_1983_Y, OR4_634_Y, OR4_2487_Y, OR4_1053_Y, OR4_2743_Y, 
        OR4_1068_Y, OR4_1347_Y, OR4_1325_Y, OR4_473_Y, OR4_1953_Y, 
        OR4_475_Y, OR4_1321_Y, OR4_318_Y, OR4_536_Y, OR4_331_Y, 
        OR4_1233_Y, OR4_2391_Y, OR4_406_Y, OR4_1811_Y, OR4_251_Y, 
        OR4_1812_Y, OR4_2660_Y, OR4_1664_Y, OR4_1883_Y, OR4_1675_Y, 
        OR4_2552_Y, OR4_708_Y, OR4_1745_Y, OR4_464_Y, OR4_1945_Y, 
        OR4_467_Y, OR4_1308_Y, OR4_303_Y, OR4_528_Y, OR4_322_Y, 
        OR4_1222_Y, OR4_2379_Y, OR2_14_Y, OR4_392_Y, OR4_1381_Y, 
        OR4_1476_Y, OR4_1372_Y, OR4_796_Y, OR4_1734_Y, OR4_2201_Y, 
        OR4_2991_Y, OR4_1858_Y, OR4_69_Y, OR4_757_Y, OR4_1083_Y, 
        OR4_2680_Y, OR4_545_Y, OR4_177_Y, OR4_1677_Y, OR4_2246_Y, 
        OR4_2079_Y, OR4_2032_Y, OR4_1069_Y, OR4_1726_Y, OR4_2038_Y, 
        OR4_601_Y, OR4_1516_Y, OR4_1188_Y, OR4_2676_Y, OR4_195_Y, 
        OR4_31_Y, OR4_3015_Y, OR4_1180_Y, OR4_1845_Y, OR4_2138_Y, 
        OR4_712_Y, OR4_1624_Y, OR4_1292_Y, OR4_2803_Y, OR4_302_Y, 
        OR4_120_Y, OR2_1_Y, OR4_2940_Y, OR4_1526_Y, OR4_1696_Y, 
        OR4_2970_Y, OR4_1552_Y, OR4_1865_Y, OR4_1689_Y, OR4_2196_Y, 
        OR4_494_Y, OR4_2604_Y, OR4_239_Y, OR4_547_Y, OR4_2139_Y, 
        OR4_36_Y, OR4_2738_Y, OR4_1193_Y, OR4_1739_Y, OR4_1563_Y, 
        OR4_1504_Y, OR4_1223_Y, OR4_1893_Y, OR4_2171_Y, OR4_751_Y, 
        OR4_1665_Y, OR4_1341_Y, OR4_2842_Y, OR4_359_Y, OR4_154_Y, 
        OR4_113_Y, OR4_1389_Y, OR4_2075_Y, OR4_2360_Y, OR4_965_Y, 
        OR4_1852_Y, OR4_1497_Y, OR4_3011_Y, OR4_541_Y, OR4_343_Y, 
        OR2_6_Y, OR4_178_Y, OR4_2471_Y, OR4_2671_Y, OR4_1013_Y, 
        OR4_327_Y, OR4_2740_Y, OR4_2212_Y, OR4_2531_Y, OR4_2990_Y, 
        OR4_2564_Y, OR4_142_Y, OR4_2371_Y, OR4_1367_Y, OR4_1641_Y, 
        OR4_1301_Y, OR4_1662_Y, OR4_2409_Y, OR4_185_Y, OR4_2281_Y, 
        OR4_1802_Y, OR4_2433_Y, OR4_1622_Y, OR4_600_Y, OR4_922_Y, 
        OR4_538_Y, OR4_953_Y, OR4_1654_Y, OR4_2475_Y, OR4_1540_Y, 
        OR4_1988_Y, OR4_2630_Y, OR4_1801_Y, OR4_774_Y, OR4_1100_Y, 
        OR4_713_Y, OR4_1118_Y, OR4_1838_Y, OR4_2674_Y, OR2_42_Y, 
        OR4_3013_Y, OR4_1892_Y, OR4_2588_Y, OR4_924_Y, OR4_1396_Y, 
        OR4_1139_Y, OR4_1170_Y, OR4_721_Y, OR4_1373_Y, OR4_2857_Y, 
        OR4_1285_Y, OR4_2861_Y, OR4_627_Y, OR4_2708_Y, OR4_2923_Y, 
        OR4_2723_Y, OR4_530_Y, OR4_1707_Y, OR4_2796_Y, OR4_1710_Y, 
        OR4_151_Y, OR4_1711_Y, OR4_2559_Y, OR4_1581_Y, OR4_1780_Y, 
        OR4_1590_Y, OR4_2457_Y, OR4_617_Y, OR4_1652_Y, OR4_2396_Y, 
        OR4_860_Y, OR4_2397_Y, OR4_193_Y, OR4_2241_Y, OR4_2461_Y, 
        OR4_2257_Y, OR4_101_Y, OR4_1310_Y, OR2_55_Y, OR4_1532_Y, 
        OR4_1853_Y, OR4_2716_Y, OR4_2773_Y, OR4_1141_Y, OR4_1307_Y, 
        OR4_194_Y, OR4_2888_Y, OR4_2997_Y, OR4_1089_Y, OR4_237_Y, 
        OR4_2194_Y, OR4_849_Y, OR4_1819_Y, OR4_2507_Y, OR4_1151_Y, 
        OR4_517_Y, OR4_2904_Y, OR4_1756_Y, OR4_1394_Y, OR4_567_Y, 
        OR4_2540_Y, OR4_1183_Y, OR4_2136_Y, OR4_2856_Y, OR4_1451_Y, 
        OR4_842_Y, OR4_147_Y, OR4_2082_Y, OR4_2204_Y, OR4_1414_Y, 
        OR4_334_Y, OR4_2005_Y, OR4_3003_Y, OR4_637_Y, OR4_2285_Y, 
        OR4_1671_Y, OR4_1032_Y, OR2_76_Y, OR4_2959_Y, OR4_696_Y, 
        OR4_2681_Y, OR4_2465_Y, OR4_2841_Y, OR4_614_Y, OR4_276_Y, 
        OR4_2045_Y, OR4_2259_Y, OR4_2795_Y, OR4_1232_Y, OR4_2798_Y, 
        OR4_564_Y, OR4_2634_Y, OR4_2858_Y, OR4_2647_Y, OR4_471_Y, 
        OR4_1642_Y, OR4_2727_Y, OR4_526_Y, OR4_2003_Y, OR4_527_Y, 
        OR4_1369_Y, OR4_377_Y, OR4_588_Y, OR4_391_Y, OR4_1274_Y, 
        OR4_2442_Y, OR4_459_Y, OR4_2497_Y, OR4_966_Y, OR4_2500_Y, 
        OR4_283_Y, OR4_2347_Y, OR4_2566_Y, OR4_2356_Y, OR4_191_Y, 
        OR4_1398_Y, OR2_60_Y, OR4_446_Y, OR4_2276_Y, OR4_867_Y, 
        OR4_222_Y, OR4_1920_Y, OR4_35_Y, OR4_384_Y, OR4_828_Y, 
        OR4_2148_Y, OR4_735_Y, OR4_300_Y, OR4_1991_Y, OR4_1426_Y, 
        OR4_2777_Y, OR4_2385_Y, OR4_409_Y, OR4_2108_Y, OR4_503_Y, 
        OR4_5_Y, OR4_2601_Y, OR4_2146_Y, OR4_789_Y, OR4_228_Y, 
        OR4_1548_Y, OR4_1217_Y, OR4_2226_Y, OR4_939_Y, OR4_2324_Y, 
        OR4_1827_Y, OR4_1166_Y, OR4_714_Y, OR4_2383_Y, OR4_1826_Y, 
        OR4_109_Y, OR4_2817_Y, OR4_813_Y, OR4_2515_Y, OR4_918_Y, 
        OR2_13_Y, OR4_2182_Y, OR4_1926_Y, OR4_1035_Y, OR4_1611_Y, 
        OR4_2918_Y, OR4_221_Y, OR4_2899_Y, OR4_855_Y, OR4_1189_Y, 
        OR4_1882_Y, OR4_2583_Y, OR4_2896_Y, OR4_1432_Y, OR4_2342_Y, 
        OR4_2001_Y, OR4_457_Y, OR4_1059_Y, OR4_861_Y, OR4_793_Y, 
        OR4_1591_Y, OR4_2274_Y, OR4_2603_Y, OR4_1173_Y, OR4_2070_Y, 
        OR4_1702_Y, OR4_158_Y, OR4_747_Y, OR4_566_Y, OR4_516_Y, 
        OR4_686_Y, OR4_1386_Y, OR4_1663_Y, OR4_234_Y, OR4_1178_Y, 
        OR4_803_Y, OR4_2287_Y, OR4_2905_Y, OR4_2711_Y, OR2_67_Y, 
        OR4_1759_Y, OR4_72_Y, OR4_1748_Y, OR4_579_Y, OR4_2145_Y, 
        OR4_805_Y, OR4_2153_Y, OR4_2445_Y, OR4_2427_Y, OR4_1438_Y, 
        OR4_2128_Y, OR4_2423_Y, OR4_1026_Y, OR4_1912_Y, OR4_1561_Y, 
        OR4_34_Y, OR4_599_Y, OR4_411_Y, OR4_355_Y, OR4_2812_Y, 
        OR4_436_Y, OR4_728_Y, OR4_2329_Y, OR4_214_Y, OR4_2933_Y, 
        OR4_1374_Y, OR4_1948_Y, OR4_1752_Y, OR4_1691_Y, OR4_1427_Y, 
        OR4_2123_Y, OR4_2414_Y, OR4_1014_Y, OR4_1904_Y, OR4_1547_Y, 
        OR4_25_Y, OR4_594_Y, OR4_398_Y, OR2_10_Y, OR4_1103_Y, 
        OR4_3034_Y, OR4_666_Y, OR4_2037_Y, OR4_2513_Y, OR4_2224_Y, 
        OR4_2261_Y, OR4_1856_Y, OR4_2482_Y, OR4_756_Y, OR4_1449_Y, 
        OR4_1744_Y, OR4_305_Y, OR4_1253_Y, OR4_897_Y, OR4_2369_Y, 
        OR4_2976_Y, OR4_2800_Y, OR4_2745_Y, OR4_2715_Y, OR4_340_Y, 
        OR4_651_Y, OR4_2231_Y, OR4_122_Y, OR4_2840_Y, OR4_1288_Y, 
        OR4_1850_Y, OR4_1657_Y, OR4_1606_Y, OR4_328_Y, OR4_1055_Y, 
        OR4_1349_Y, OR4_2956_Y, OR4_812_Y, OR4_458_Y, OR4_1957_Y, 
        OR4_2535_Y, OR4_2337_Y, OR2_53_Y, OR4_2577_Y, OR4_1155_Y, 
        OR4_2085_Y, OR4_1757_Y, OR4_2219_Y, OR4_163_Y, OR4_2240_Y, 
        OR4_762_Y, OR4_1357_Y, OR4_2389_Y, OR4_847_Y, OR4_2390_Y, 
        OR4_181_Y, OR4_2235_Y, OR4_2455_Y, OR4_2245_Y, OR4_90_Y, 
        OR4_1300_Y, OR4_2320_Y, OR4_993_Y, OR4_2441_Y, OR4_996_Y, 
        OR4_1797_Y, OR4_830_Y, OR4_1056_Y, OR4_850_Y, OR4_1697_Y, 
        OR4_2930_Y, OR4_926_Y, OR4_1922_Y, OR4_357_Y, OR4_1924_Y, 
        OR4_2781_Y, OR4_1768_Y, OR4_1981_Y, OR4_1779_Y, OR4_2672_Y, 
        OR4_810_Y, OR2_45_Y, OR4_2821_Y, OR4_2087_Y, OR4_1500_Y, 
        OR4_1935_Y, OR4_1866_Y, OR4_116_Y, OR4_2898_Y, OR4_452_Y, 
        OR4_1934_Y, OR4_2126_Y, OR4_2793_Y, OR4_1954_Y, OR4_954_Y, 
        OR4_1245_Y, OR4_879_Y, OR4_1261_Y, OR4_1989_Y, OR4_2829_Y, 
        OR4_1867_Y, OR4_1418_Y, OR4_2053_Y, OR4_1255_Y, OR4_200_Y, 
        OR4_518_Y, OR4_133_Y, OR4_531_Y, OR4_1291_Y, OR4_2092_Y, 
        OR4_1172_Y, OR4_843_Y, OR4_1462_Y, OR4_663_Y, OR4_2684_Y, 
        OR4_2984_Y, OR4_2613_Y, OR4_2998_Y, OR4_700_Y, OR4_1502_Y, 
        OR2_15_Y, OR4_388_Y, OR4_2345_Y, OR4_783_Y, OR4_281_Y, 
        OR4_1979_Y, OR4_81_Y, OR4_444_Y, OR4_753_Y, OR4_2203_Y, 
        OR4_683_Y, OR4_245_Y, OR4_1932_Y, OR4_1378_Y, OR4_2706_Y, 
        OR4_2317_Y, OR4_337_Y, OR4_2050_Y, OR4_427_Y, OR4_2981_Y, 
        OR4_2658_Y, OR4_2197_Y, OR4_872_Y, OR4_288_Y, OR4_1610_Y, 
        OR4_1272_Y, OR4_2301_Y, OR4_1003_Y, OR4_2394_Y, OR4_1897_Y, 
        OR4_1102_Y, OR4_662_Y, OR4_2315_Y, OR4_1762_Y, OR4_56_Y, 
        OR4_2758_Y, OR4_739_Y, OR4_2444_Y, OR4_845_Y, OR2_8_Y, 
        OR4_2511_Y, OR4_1162_Y, OR4_1054_Y, OR4_2616_Y, OR4_1863_Y, 
        OR4_2897_Y, OR4_2325_Y, OR4_2726_Y, OR4_2774_Y, OR4_2831_Y, 
        OR4_2365_Y, OR4_1040_Y, OR4_451_Y, OR4_1766_Y, OR4_1417_Y, 
        OR4_2464_Y, OR4_1153_Y, OR4_2561_Y, OR4_2057_Y, OR4_1437_Y, 
        OR4_1037_Y, OR4_2702_Y, OR4_2121_Y, OR4_405_Y, OR4_54_Y, 
        OR4_1121_Y, OR4_2833_Y, OR4_1212_Y, OR4_691_Y, OR4_1344_Y, 
        OR4_912_Y, OR4_2582_Y, OR4_2016_Y, OR4_284_Y, OR4_2989_Y, 
        OR4_1015_Y, OR4_2712_Y, OR4_1097_Y, OR2_16_Y, OR4_811_Y, 
        OR4_1512_Y, OR4_1284_Y, OR4_557_Y, OR4_646_Y, OR4_2501_Y, 
        OR4_2040_Y, OR4_1107_Y, OR4_1740_Y, OR4_332_Y, OR4_2570_Y, 
        OR4_1490_Y, OR4_111_Y, OR4_1120_Y, OR4_1778_Y, OR4_413_Y, 
        OR4_2853_Y, OR4_2144_Y, OR4_1061_Y, OR4_1067_Y, OR4_218_Y, 
        OR4_2176_Y, OR4_822_Y, OR4_1799_Y, OR4_2479_Y, OR4_1134_Y, 
        OR4_496_Y, OR4_2874_Y, OR4_1725_Y, OR4_802_Y, OR4_3037_Y, 
        OR4_1960_Y, OR4_577_Y, OR4_1566_Y, OR4_2223_Y, OR4_890_Y, 
        OR4_244_Y, OR4_2623_Y, OR2_36_Y, OR4_1050_Y, OR4_1810_Y, 
        OR4_745_Y, OR4_560_Y, OR4_923_Y, OR4_1727_Y, OR4_1411_Y, 
        OR4_127_Y, OR4_362_Y, OR4_702_Y, OR4_1401_Y, OR4_1681_Y, 
        OR4_248_Y, OR4_1196_Y, OR4_827_Y, OR4_2303_Y, OR4_2926_Y, 
        OR4_2731_Y, OR4_2667_Y, OR4_1483_Y, OR4_2167_Y, OR4_2477_Y, 
        OR4_1071_Y, OR4_1965_Y, OR4_1607_Y, OR4_70_Y, OR4_654_Y, 
        OR4_465_Y, OR4_407_Y, OR4_422_Y, OR4_1140_Y, OR4_1420_Y, 
        OR4_3038_Y, OR4_919_Y, OR4_553_Y, OR4_2046_Y, OR4_2635_Y, 
        OR4_2429_Y, OR2_57_Y, OR4_2547_Y, OR4_24_Y, OR4_2217_Y, 
        OR4_58_Y, OR4_1000_Y, OR4_1928_Y, OR4_1094_Y, OR4_1412_Y, 
        OR4_3020_Y, OR4_1881_Y, OR4_2512_Y, OR4_1686_Y, OR4_673_Y, 
        OR4_999_Y, OR4_604_Y, OR4_1016_Y, OR4_1720_Y, OR4_2548_Y, 
        OR4_1605_Y, OR4_2366_Y, OR4_3029_Y, OR4_2177_Y, OR4_1195_Y, 
        OR4_1465_Y, OR4_1123_Y, OR4_1484_Y, OR4_2207_Y, OR4_27_Y, 
        OR4_2107_Y, OR4_1578_Y, OR4_2188_Y, OR4_1403_Y, OR4_365_Y, 
        OR4_672_Y, OR4_292_Y, OR4_692_Y, OR4_1429_Y, OR4_2222_Y, 
        OR2_31_Y, OR4_2025_Y, OR4_1445_Y, OR4_1186_Y, OR4_2682_Y, 
        OR4_607_Y, OR4_2307_Y, OR4_1213_Y, OR4_1402_Y, OR4_1029_Y, 
        OR4_1849_Y, OR4_285_Y, OR4_1854_Y, OR4_2705_Y, OR4_1698_Y, 
        OR4_1917_Y, OR4_1708_Y, OR4_2605_Y, OR4_734_Y, OR4_1783_Y, 
        OR4_1294_Y, OR4_2789_Y, OR4_1296_Y, OR4_2110_Y, OR4_1157_Y, 
        OR4_1359_Y, OR4_1171_Y, OR4_2023_Y, OR4_157_Y, OR4_1242_Y, 
        OR4_1023_Y, OR4_2470_Y, OR4_1027_Y, OR4_1823_Y, OR4_871_Y, 
        OR4_1081_Y, OR4_881_Y, OR4_1722_Y, OR4_2945_Y, OR2_29_Y, 
        OR4_1163_Y, OR4_831_Y, OR4_690_Y, OR4_2865_Y, OR4_311_Y, 
        OR4_1278_Y, OR4_77_Y, OR4_2159_Y, OR4_1985_Y, OR4_479_Y, 
        OR4_1131_Y, OR4_291_Y, OR4_2295_Y, OR4_2619_Y, OR4_2218_Y, 
        OR4_2638_Y, OR4_326_Y, OR4_1168_Y, OR4_199_Y, OR4_145_Y, 
        OR4_790_Y, OR4_3032_Y, OR4_1992_Y, OR4_2280_Y, OR4_1929_Y, 
        OR4_2298_Y, OR4_32_Y, OR4_836_Y, OR4_2954_Y, OR4_33_Y, 
        OR4_657_Y, OR4_2902_Y, OR4_1843_Y, OR4_2142_Y, OR4_1774_Y, 
        OR4_2152_Y, OR4_2939_Y, OR4_698_Y, OR2_71_Y, OR4_2752_Y, 
        OR4_877_Y, OR4_2609_Y, OR4_1430_Y, OR4_2272_Y, OR4_1513_Y, 
        OR4_1279_Y, OR4_763_Y, OR4_737_Y, OR4_2556_Y, OR4_1028_Y, 
        OR4_2558_Y, OR4_346_Y, OR4_2403_Y, OR4_2627_Y, OR4_2417_Y, 
        OR4_252_Y, OR4_1444_Y, OR4_2494_Y, OR4_697_Y, OR4_2154_Y, 
        OR4_699_Y, OR4_1523_Y, OR4_552_Y, OR4_746_Y, OR4_561_Y, 
        OR4_1424_Y, OR4_2624_Y, OR4_629_Y, OR4_2420_Y, OR4_887_Y, 
        OR4_2421_Y, OR4_220_Y, OR4_2269_Y, OR4_2490_Y, OR4_2286_Y, 
        OR4_124_Y, OR4_1335_Y, OR2_56_Y, OR4_511_Y, OR4_1909_Y, 
        OR4_2975_Y, OR4_2808_Y, OR4_1425_Y, OR4_182_Y, OR4_2881_Y, 
        OR4_1289_Y, OR4_533_Y, OR4_48_Y, OR4_2236_Y, OR4_1211_Y, 
        OR4_2869_Y, OR4_798_Y, OR4_1477_Y, OR4_106_Y, OR4_2530_Y, 
        OR4_1847_Y, OR4_724_Y, OR4_1436_Y, OR4_622_Y, OR4_2608_Y, 
        OR4_1238_Y, OR4_2181_Y, OR4_2910_Y, OR4_1511_Y, OR4_905_Y, 
        OR4_209_Y, OR4_2129_Y, OR4_2485_Y, OR4_1659_Y, OR4_608_Y, 
        OR4_2242_Y, OR4_204_Y, OR4_910_Y, OR4_2567_Y, OR4_1943_Y, 
        OR4_1280_Y, OR2_4_Y, OR4_1715_Y, OR4_740_Y, OR4_609_Y, 
        OR4_383_Y, OR4_238_Y, OR4_1841_Y, OR4_14_Y, OR4_2786_Y, 
        OR4_1908_Y, OR4_1562_Y, OR4_19_Y, OR4_1564_Y, OR4_2387_Y, 
        OR4_1419_Y, OR4_1618_Y, OR4_1428_Y, OR4_2288_Y, OR4_448_Y, 
        OR4_1492_Y, OR4_582_Y, OR4_2066_Y, OR4_584_Y, OR4_1416_Y, 
        OR4_431_Y, OR4_648_Y, OR4_447_Y, OR4_1336_Y, OR4_2509_Y, 
        OR4_524_Y, OR4_432_Y, OR4_1923_Y, OR4_435_Y, OR4_1290_Y, 
        OR4_290_Y, OR4_509_Y, OR4_295_Y, OR4_1199_Y, OR4_2358_Y, 
        OR2_12_Y, OR4_661_Y, OR4_2243_Y, OR4_159_Y, OR4_2915_Y, 
        OR4_324_Y, OR4_1322_Y, OR4_341_Y, OR4_1894_Y, OR4_2462_Y, 
        OR4_316_Y, OR4_1047_Y, OR4_1334_Y, OR4_2943_Y, OR4_799_Y, 
        OR4_445_Y, OR4_1949_Y, OR4_2528_Y, OR4_2323_Y, OR4_2267_Y, 
        OR4_1941_Y, OR4_2644_Y, OR4_2952_Y, OR4_1489_Y, OR4_2399_Y, 
        OR4_2065_Y, OR4_523_Y, OR4_1114_Y, OR4_931_Y, OR4_874_Y, 
        OR4_2916_Y, OR4_546_Y, OR4_853_Y, OR4_2436_Y, OR4_310_Y, 
        OR4_3024_Y, OR4_1459_Y, OR4_2047_Y, OR4_1859_Y, OR2_44_Y, 
        OR4_2901_Y, OR4_2767_Y, OR4_1913_Y, OR4_2536_Y, OR4_2571_Y, 
        OR4_1574_Y, OR4_2524_Y, OR4_701_Y, OR4_1022_Y, OR4_2729_Y, 
        OR4_1164_Y, OR4_2730_Y, OR4_507_Y, OR4_2573_Y, OR4_2797_Y, 
        OR4_2589_Y, OR4_404_Y, OR4_1592_Y, OR4_2653_Y, OR4_2594_Y, 
        OR4_1042_Y, OR4_2595_Y, OR4_370_Y, OR4_2425_Y, OR4_2651_Y, 
        OR4_2437_Y, OR4_272_Y, OR4_1460_Y, OR4_2514_Y, OR4_1733_Y, 
        OR4_172_Y, OR4_1736_Y, OR4_2596_Y, OR4_1598_Y, OR4_1805_Y, 
        OR4_1609_Y, OR4_2478_Y, OR4_640_Y, OR2_41_Y, OR4_2056_Y, 
        OR4_2_Y, OR4_98_Y, OR4_3035_Y, OR4_2451_Y, OR4_363_Y, 
        OR4_857_Y, OR4_1594_Y, OR4_482_Y, OR4_1393_Y, OR4_2022_Y, 
        OR4_1228_Y, OR4_164_Y, OR4_485_Y, OR4_108_Y, OR4_505_Y, 
        OR4_1257_Y, OR4_2061_Y, OR4_1138_Y, OR4_2352_Y, OR4_3007_Y, 
        OR4_2161_Y, OR4_1176_Y, OR4_1450_Y, OR4_1105_Y, OR4_1464_Y, 
        OR4_2192_Y, OR4_10_Y, OR4_2094_Y, OR4_2467_Y, OR4_68_Y, 
        OR4_2279_Y, OR4_1281_Y, OR4_1570_Y, OR4_1224_Y, OR4_1582_Y, 
        OR4_2314_Y, OR4_102_Y, OR2_50_Y, OR4_1535_Y, OR4_136_Y, 
        OR4_314_Y, OR4_1572_Y, OR4_160_Y, OR4_490_Y, OR4_306_Y, 
        OR4_851_Y, OR4_2140_Y, OR4_886_Y, OR4_1498_Y, OR4_694_Y, 
        OR4_2722_Y, OR4_3018_Y, OR4_2645_Y, OR4_3036_Y, OR4_718_Y, 
        OR4_1538_Y, OR4_602_Y, OR4_2517_Y, OR4_107_Y, OR4_2322_Y, 
        OR4_1328_Y, OR4_1608_Y, OR4_1262_Y, OR4_1623_Y, OR4_2362_Y, 
        OR4_138_Y, OR4_2229_Y, OR4_2717_Y, OR4_282_Y, OR4_2516_Y, 
        OR4_1482_Y, OR4_1786_Y, OR4_1423_Y, OR4_1806_Y, OR4_2551_Y, 
        OR4_320_Y, OR2_59_Y, OR4_2835_Y, OR4_2868_Y, OR4_55_Y, 
        OR4_1626_Y, OR4_1388_Y, OR4_2258_Y, OR4_4_Y, OR4_1518_Y, 
        OR4_2341_Y, OR4_2331_Y, OR4_1524_Y, OR4_461_Y, OR4_2114_Y, 
        OR4_66_Y, OR4_743_Y, OR4_2402_Y, OR4_1787_Y, OR4_1136_Y, 
        OR4_17_Y, OR4_2364_Y, OR4_1557_Y, OR4_499_Y, OR4_2141_Y, 
        OR4_96_Y, OR4_778_Y, OR4_2440_Y, OR4_1820_Y, OR4_1175_Y, 
        OR4_46_Y, OR4_2626_Y, OR4_1793_Y, OR4_726_Y, OR4_2388_Y, 
        OR4_335_Y, OR4_1051_Y, OR4_2710_Y, OR4_2072_Y, OR4_1405_Y, 
        OR2_5_Y, CFG3_17_Y, CFG3_5_Y, CFG3_10_Y, CFG3_23_Y, CFG3_4_Y, 
        CFG3_1_Y, CFG3_0_Y, CFG3_13_Y, CFG3_14_Y, CFG3_7_Y, CFG3_3_Y, 
        CFG3_18_Y, OR4_105_Y, OR4_2593_Y, OR4_2277_Y, OR4_748_Y, 
        OR4_1717_Y, OR4_408_Y, OR4_2306_Y, OR4_2523_Y, OR4_2124_Y, 
        OR4_2845_Y, OR4_481_Y, OR4_769_Y, OR4_2370_Y, OR4_249_Y, 
        OR4_2965_Y, OR4_1409_Y, OR4_1980_Y, OR4_1788_Y, OR4_1728_Y, 
        OR4_2230_Y, OR4_2967_Y, OR4_196_Y, OR4_1803_Y, OR4_2750_Y, 
        OR4_2361_Y, OR4_834_Y, OR4_1415_Y, OR4_1243_Y, OR4_1192_Y, 
        OR4_1966_Y, OR4_2675_Y, OR4_2973_Y, OR4_1522_Y, OR4_2432_Y, 
        OR4_2086_Y, OR4_548_Y, OR4_1145_Y, OR4_962_Y, OR2_26_Y, 
        OR4_652_Y, OR4_168_Y, OR4_1295_Y, OR4_1259_Y, OR4_2932_Y, 
        OR4_839_Y, OR4_114_Y, OR4_2880_Y, OR4_983_Y, OR4_167_Y, 
        OR4_2393_Y, OR4_1354_Y, OR4_3005_Y, OR4_971_Y, OR4_1619_Y, 
        OR4_243_Y, OR4_2685_Y, OR4_1997_Y, OR4_894_Y, OR4_2779_Y, 
        OR4_1937_Y, OR4_884_Y, OR4_2529_Y, OR4_477_Y, OR4_1181_Y, 
        OR4_2846_Y, OR4_2179_Y, OR4_1527_Y, OR4_410_Y, OR4_816_Y, 
        OR4_12_Y, OR4_1969_Y, OR4_591_Y, OR4_1579_Y, OR4_2237_Y, 
        OR4_900_Y, OR4_260_Y, OR4_2637_Y, OR2_37_Y, OR4_2084_Y, 
        OR4_2299_Y, OR4_71_Y, OR4_899_Y, OR4_960_Y, OR4_395_Y, 
        OR4_1545_Y, OR4_1712_Y, OR4_2791_Y, OR4_1916_Y, OR4_354_Y, 
        OR4_1921_Y, OR4_2776_Y, OR4_1765_Y, OR4_1977_Y, OR4_1777_Y, 
        OR4_2668_Y, OR4_807_Y, OR4_1851_Y, OR4_2134_Y, OR4_586_Y, 
        OR4_2135_Y, OR4_2993_Y, OR4_2002_Y, OR4_2186_Y, OR4_2018_Y, 
        OR4_2907_Y, OR4_1057_Y, OR4_2080_Y, OR4_2961_Y, OR4_1391_Y, 
        OR4_2963_Y, OR4_725_Y, OR4_2818_Y, OR4_3019_Y, OR4_2834_Y, 
        OR4_645_Y, OR4_1824_Y, OR2_74_Y, OR4_1546_Y, OR4_2200_Y, 
        OR4_2228_Y, OR4_2669_Y, OR4_2198_Y, OR4_250_Y, OR4_1844_Y, 
        OR4_2248_Y, OR4_650_Y, OR4_1099_Y, OR4_261_Y, OR4_2213_Y, 
        OR4_875_Y, OR4_1839_Y, OR4_2532_Y, OR4_1174_Y, OR4_532_Y, 
        OR4_2927_Y, OR4_1770_Y, OR4_1749_Y, OR4_964_Y, OR4_2937_Y, 
        OR4_1530_Y, OR4_2521_Y, OR4_149_Y, OR4_1821_Y, OR4_1229_Y, 
        OR4_534_Y, OR4_2446_Y, OR4_1773_Y, OR4_985_Y, OR4_2960_Y, 
        OR4_1554_Y, OR4_2545_Y, OR4_174_Y, OR4_1848_Y, OR4_1248_Y, 
        OR4_559_Y, OR2_62_Y, OR4_7_Y, OR4_2599_Y, OR4_908_Y, 
        OR4_2928_Y, OR4_1661_Y, OR4_1961_Y, OR4_1431_Y, OR4_2526_Y, 
        OR4_345_Y, OR4_2885_Y, OR4_1320_Y, OR4_2889_Y, OR4_664_Y, 
        OR4_2746_Y, OR4_2948_Y, OR4_2757_Y, OR4_565_Y, OR4_1746_Y, 
        OR4_2822_Y, OR4_2405_Y, OR4_873_Y, OR4_2408_Y, OR4_198_Y, 
        OR4_2254_Y, OR4_2474_Y, OR4_2268_Y, OR4_110_Y, OR4_1324_Y, 
        OR4_2344_Y, OR4_717_Y, OR4_2184_Y, OR4_720_Y, OR4_1556_Y, 
        OR4_583_Y, OR4_781_Y, OR4_595_Y, OR4_1455_Y, OR4_2664_Y, 
        OR2_20_Y, OR4_817_Y, OR4_1984_Y, OR4_689_Y, OR4_2560_Y, 
        OR4_373_Y, OR4_2649_Y, OR4_2381_Y, OR4_1896_Y, OR4_1874_Y, 
        OR4_492_Y, OR4_1204_Y, OR4_1472_Y, OR4_51_Y, OR4_981_Y, 
        OR4_610_Y, OR4_2098_Y, OR4_2703_Y, OR4_2498_Y, OR4_2435_Y, 
        OR4_1645_Y, OR4_2346_Y, OR4_2661_Y, OR4_1240_Y, OR4_2127_Y, 
        OR4_1771_Y, OR4_233_Y, OR4_825_Y, OR4_635_Y, OR4_574_Y, 
        OR4_358_Y, OR4_1075_Y, OR4_1366_Y, OR4_2972_Y, OR4_837_Y, 
        OR4_484_Y, OR4_1973_Y, OR4_2555_Y, OR4_2359_Y, OR2_54_Y, 
        OR4_2051_Y, OR4_1286_Y, OR4_2867_Y, OR4_927_Y, OR4_906_Y, 
        OR4_86_Y, OR4_2575_Y, OR4_2027_Y, OR4_1148_Y, OR4_2334_Y, 
        OR4_1915_Y, OR4_556_Y, OR4_3_Y, OR4_1329_Y, OR4_978_Y, 
        OR4_2012_Y, OR4_677_Y, OR4_2095_Y, OR4_1586_Y, OR4_1569_Y, 
        OR4_1156_Y, OR4_2836_Y, OR4_2233_Y, OR4_537_Y, OR4_162_Y, 
        OR4_1249_Y, OR4_2958_Y, OR4_1339_Y, OR4_819_Y, OR4_94_Y, 
        OR4_2736_Y, OR4_1361_Y, OR4_780_Y, OR4_2100_Y, OR4_1738_Y, 
        OR4_2827_Y, OR4_1461_Y, OR4_2920_Y, OR2_58_Y, OR4_2872_Y, 
        OR4_1878_Y, OR4_1721_Y, OR4_1510_Y, OR4_1382_Y, OR4_2988_Y, 
        OR4_1142_Y, OR4_859_Y, OR4_13_Y, OR4_2534_Y, OR4_171_Y, 
        OR4_487_Y, OR4_2088_Y, OR4_3017_Y, OR4_2662_Y, OR4_1126_Y, 
        OR4_1680_Y, OR4_1496_Y, OR4_1443_Y, OR4_1544_Y, OR4_2221_Y, 
        OR4_2542_Y, OR4_1124_Y, OR4_2028_Y, OR4_1660_Y, OR4_123_Y, 
        OR4_709_Y, OR4_525_Y, OR4_470_Y, OR4_1413_Y, OR4_2096_Y, 
        OR4_2392_Y, OR4_991_Y, OR4_1886_Y, OR4_1529_Y, OR4_0_Y, 
        OR4_568_Y, OR4_379_Y, OR2_7_Y, OR4_982_Y, OR4_838_Y, OR4_18_Y, 
        OR4_624_Y, OR4_653_Y, OR4_2719_Y, OR4_612_Y, OR4_1816_Y, 
        OR4_2117_Y, OR4_639_Y, OR4_1350_Y, OR4_1621_Y, OR4_183_Y, 
        OR4_1128_Y, OR4_749_Y, OR4_2234_Y, OR4_2862_Y, OR4_2657_Y, 
        OR4_2606_Y, OR4_512_Y, OR4_1227_Y, OR4_1493_Y, OR4_64_Y, 
        OR4_1008_Y, OR4_633_Y, OR4_2122_Y, OR4_2728_Y, OR4_2518_Y, 
        OR4_2458_Y, OR4_2742_Y, OR4_367_Y, OR4_671_Y, OR4_2252_Y, 
        OR4_137_Y, OR4_2863_Y, OR4_1305_Y, OR4_1876_Y, OR4_1674_Y, 
        OR2_40_Y, OR4_829_Y, OR4_543_Y, OR4_2683_Y, OR4_232_Y, 
        OR4_1508_Y, OR4_1890_Y, OR4_1486_Y, OR4_2505_Y, OR4_2850_Y, 
        OR4_141_Y, OR4_784_Y, OR4_3031_Y, OR4_1987_Y, OR4_2275_Y, 
        OR4_1927_Y, OR4_2294_Y, OR4_26_Y, OR4_832_Y, OR4_2949_Y, 
        OR4_2938_Y, OR4_510_Y, OR4_2755_Y, OR4_1694_Y, OR4_2009_Y, 
        OR4_1628_Y, OR4_2030_Y, OR4_2794_Y, OR4_549_Y, OR4_2656_Y, 
        OR4_2000_Y, OR4_2643_Y, OR4_1813_Y, OR4_786_Y, OR4_1112_Y, 
        OR4_719_Y, OR4_1133_Y, OR4_1855_Y, OR4_2687_Y, OR2_43_Y, 
        OR4_387_Y, OR4_1716_Y, OR4_374_Y, OR4_2214_Y, OR4_771_Y, 
        OR4_2460_Y, OR4_785_Y, OR4_1095_Y, OR4_1079_Y, OR4_2785_Y, 
        OR4_344_Y, OR4_2592_Y, OR4_1542_Y, OR4_1846_Y, OR4_1479_Y, 
        OR4_1870_Y, OR4_2620_Y, OR4_390_Y, OR4_2488_Y, OR4_1088_Y, 
        OR4_1685_Y, OR4_898_Y, OR4_2924_Y, OR4_146_Y, OR4_2854_Y, 
        OR4_161_Y, OR4_949_Y, OR4_1723_Y, OR4_795_Y, OR4_2769_Y, 
        OR4_333_Y, OR4_2578_Y, OR4_1537_Y, OR4_1837_Y, OR4_1467_Y, 
        OR4_1860_Y, OR4_2614_Y, OR4_380_Y, OR2_63_Y, OR4_2770_Y, 
        OR4_1629_Y, OR4_2309_Y, OR4_660_Y, OR4_1150_Y, OR4_885_Y, 
        OR4_914_Y, OR4_478_Y, OR4_1127_Y, OR4_2077_Y, OR4_2737_Y, 
        OR4_1901_Y, OR4_888_Y, OR4_1197_Y, OR4_806_Y, OR4_1207_Y, 
        OR4_1938_Y, OR4_2778_Y, OR4_1807_Y, OR4_997_Y, OR4_1602_Y, 
        OR4_787_Y, OR4_2826_Y, OR4_67_Y, OR4_2760_Y, OR4_82_Y, 
        OR4_833_Y, OR4_1633_Y, OR4_706_Y, OR4_1639_Y, OR4_2271_Y, 
        OR4_1463_Y, OR4_441_Y, OR4_742_Y, OR4_381_Y, OR4_759_Y, 
        OR4_1506_Y, OR4_2310_Y, OR2_32_Y, VCC, GND, ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    OR4 OR4_1629 (.A(OR4_1127_Y), .B(OR4_2077_Y), .C(OR4_2737_Y), .D(
        OR4_1901_Y), .Y(OR4_1629_Y));
    OR4 OR4_1532 (.A(OR4_1141_Y), .B(OR4_1307_Y), .C(OR4_194_Y), .D(
        OR4_2888_Y), .Y(OR4_1532_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%82%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R82C2 (
        .A_DOUT({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, 
        nc10, nc11, nc12, nc13, nc14, \A_DOUT_TEMPR82[14] , 
        \A_DOUT_TEMPR82[13] , \A_DOUT_TEMPR82[12] , 
        \A_DOUT_TEMPR82[11] , \A_DOUT_TEMPR82[10] }), .B_DOUT({nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27, nc28, nc29, \B_DOUT_TEMPR82[14] , 
        \B_DOUT_TEMPR82[13] , \B_DOUT_TEMPR82[12] , 
        \B_DOUT_TEMPR82[11] , \B_DOUT_TEMPR82[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[82][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_387 (.A(OR4_771_Y), .B(OR4_2460_Y), .C(OR4_785_Y), .D(
        OR4_1095_Y), .Y(OR4_387_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%9%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R9C4 (
        .A_DOUT({nc30, nc31, nc32, nc33, nc34, nc35, nc36, nc37, nc38, 
        nc39, nc40, nc41, nc42, nc43, nc44, \A_DOUT_TEMPR9[24] , 
        \A_DOUT_TEMPR9[23] , \A_DOUT_TEMPR9[22] , \A_DOUT_TEMPR9[21] , 
        \A_DOUT_TEMPR9[20] }), .B_DOUT({nc45, nc46, nc47, nc48, nc49, 
        nc50, nc51, nc52, nc53, nc54, nc55, nc56, nc57, nc58, nc59, 
        \B_DOUT_TEMPR9[24] , \B_DOUT_TEMPR9[23] , \B_DOUT_TEMPR9[22] , 
        \B_DOUT_TEMPR9[21] , \B_DOUT_TEMPR9[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[9][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_888 (.A(\B_DOUT_TEMPR87[26] ), .B(\B_DOUT_TEMPR88[26] ), 
        .C(\B_DOUT_TEMPR89[26] ), .D(\B_DOUT_TEMPR90[26] ), .Y(
        OR4_888_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%94%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R94C3 (
        .A_DOUT({nc60, nc61, nc62, nc63, nc64, nc65, nc66, nc67, nc68, 
        nc69, nc70, nc71, nc72, nc73, nc74, \A_DOUT_TEMPR94[19] , 
        \A_DOUT_TEMPR94[18] , \A_DOUT_TEMPR94[17] , 
        \A_DOUT_TEMPR94[16] , \A_DOUT_TEMPR94[15] }), .B_DOUT({nc75, 
        nc76, nc77, nc78, nc79, nc80, nc81, nc82, nc83, nc84, nc85, 
        nc86, nc87, nc88, nc89, \B_DOUT_TEMPR94[19] , 
        \B_DOUT_TEMPR94[18] , \B_DOUT_TEMPR94[17] , 
        \B_DOUT_TEMPR94[16] , \B_DOUT_TEMPR94[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[94][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1182 (.A(\A_DOUT_TEMPR24[27] ), .B(\A_DOUT_TEMPR25[27] ), 
        .C(\A_DOUT_TEMPR26[27] ), .D(\A_DOUT_TEMPR27[27] ), .Y(
        OR4_1182_Y));
    OR4 OR4_681 (.A(\A_DOUT_TEMPR95[25] ), .B(\A_DOUT_TEMPR96[25] ), 
        .C(\A_DOUT_TEMPR97[25] ), .D(\A_DOUT_TEMPR98[25] ), .Y(
        OR4_681_Y));
    OR4 OR4_2355 (.A(OR4_400_Y), .B(OR4_208_Y), .C(OR4_148_Y), .D(
        OR4_495_Y), .Y(OR4_2355_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%6%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R6C5 (
        .A_DOUT({nc90, nc91, nc92, nc93, nc94, nc95, nc96, nc97, nc98, 
        nc99, nc100, nc101, nc102, nc103, nc104, \A_DOUT_TEMPR6[29] , 
        \A_DOUT_TEMPR6[28] , \A_DOUT_TEMPR6[27] , \A_DOUT_TEMPR6[26] , 
        \A_DOUT_TEMPR6[25] }), .B_DOUT({nc105, nc106, nc107, nc108, 
        nc109, nc110, nc111, nc112, nc113, nc114, nc115, nc116, nc117, 
        nc118, nc119, \B_DOUT_TEMPR6[29] , \B_DOUT_TEMPR6[28] , 
        \B_DOUT_TEMPR6[27] , \B_DOUT_TEMPR6[26] , \B_DOUT_TEMPR6[25] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[6][5] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[29], A_DIN[28], A_DIN[27], 
        A_DIN[26], A_DIN[25]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2918 (.A(OR4_2274_Y), .B(OR4_2603_Y), .C(OR4_1173_Y), .D(
        OR4_2070_Y), .Y(OR4_2918_Y));
    OR4 OR4_699 (.A(\B_DOUT_TEMPR4[18] ), .B(\B_DOUT_TEMPR5[18] ), .C(
        \B_DOUT_TEMPR6[18] ), .D(\B_DOUT_TEMPR7[18] ), .Y(OR4_699_Y));
    OR4 \OR4_B_DOUT[2]  (.A(OR4_1546_Y), .B(OR4_2200_Y), .C(OR4_2228_Y)
        , .D(OR4_2669_Y), .Y(B_DOUT[2]));
    OR4 OR4_215 (.A(\A_DOUT_TEMPR24[33] ), .B(\A_DOUT_TEMPR25[33] ), 
        .C(\A_DOUT_TEMPR26[33] ), .D(\A_DOUT_TEMPR27[33] ), .Y(
        OR4_215_Y));
    OR4 \OR4_A_DOUT[4]  (.A(OR4_2051_Y), .B(OR4_1286_Y), .C(OR4_2867_Y)
        , .D(OR4_927_Y), .Y(A_DOUT[4]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%50%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R50C0 (
        .A_DOUT({nc120, nc121, nc122, nc123, nc124, nc125, nc126, 
        nc127, nc128, nc129, nc130, nc131, nc132, nc133, nc134, 
        \A_DOUT_TEMPR50[4] , \A_DOUT_TEMPR50[3] , \A_DOUT_TEMPR50[2] , 
        \A_DOUT_TEMPR50[1] , \A_DOUT_TEMPR50[0] }), .B_DOUT({nc135, 
        nc136, nc137, nc138, nc139, nc140, nc141, nc142, nc143, nc144, 
        nc145, nc146, nc147, nc148, nc149, \B_DOUT_TEMPR50[4] , 
        \B_DOUT_TEMPR50[3] , \B_DOUT_TEMPR50[2] , \B_DOUT_TEMPR50[1] , 
        \B_DOUT_TEMPR50[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%55%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R55C4 (
        .A_DOUT({nc150, nc151, nc152, nc153, nc154, nc155, nc156, 
        nc157, nc158, nc159, nc160, nc161, nc162, nc163, nc164, 
        \A_DOUT_TEMPR55[24] , \A_DOUT_TEMPR55[23] , 
        \A_DOUT_TEMPR55[22] , \A_DOUT_TEMPR55[21] , 
        \A_DOUT_TEMPR55[20] }), .B_DOUT({nc165, nc166, nc167, nc168, 
        nc169, nc170, nc171, nc172, nc173, nc174, nc175, nc176, nc177, 
        nc178, nc179, \B_DOUT_TEMPR55[24] , \B_DOUT_TEMPR55[23] , 
        \B_DOUT_TEMPR55[22] , \B_DOUT_TEMPR55[21] , 
        \B_DOUT_TEMPR55[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[55][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_76 (.A(\B_DOUT_TEMPR72[1] ), .B(\B_DOUT_TEMPR73[1] ), .Y(
        OR2_76_Y));
    OR4 OR4_48 (.A(\B_DOUT_TEMPR75[0] ), .B(\B_DOUT_TEMPR76[0] ), .C(
        \B_DOUT_TEMPR77[0] ), .D(\B_DOUT_TEMPR78[0] ), .Y(OR4_48_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%83%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R83C1 (
        .A_DOUT({nc180, nc181, nc182, nc183, nc184, nc185, nc186, 
        nc187, nc188, nc189, nc190, nc191, nc192, nc193, nc194, 
        \A_DOUT_TEMPR83[9] , \A_DOUT_TEMPR83[8] , \A_DOUT_TEMPR83[7] , 
        \A_DOUT_TEMPR83[6] , \A_DOUT_TEMPR83[5] }), .B_DOUT({nc195, 
        nc196, nc197, nc198, nc199, nc200, nc201, nc202, nc203, nc204, 
        nc205, nc206, nc207, nc208, nc209, \B_DOUT_TEMPR83[9] , 
        \B_DOUT_TEMPR83[8] , \B_DOUT_TEMPR83[7] , \B_DOUT_TEMPR83[6] , 
        \B_DOUT_TEMPR83[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[83][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%24%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R24C2 (
        .A_DOUT({nc210, nc211, nc212, nc213, nc214, nc215, nc216, 
        nc217, nc218, nc219, nc220, nc221, nc222, nc223, nc224, 
        \A_DOUT_TEMPR24[14] , \A_DOUT_TEMPR24[13] , 
        \A_DOUT_TEMPR24[12] , \A_DOUT_TEMPR24[11] , 
        \A_DOUT_TEMPR24[10] }), .B_DOUT({nc225, nc226, nc227, nc228, 
        nc229, nc230, nc231, nc232, nc233, nc234, nc235, nc236, nc237, 
        nc238, nc239, \B_DOUT_TEMPR24[14] , \B_DOUT_TEMPR24[13] , 
        \B_DOUT_TEMPR24[12] , \B_DOUT_TEMPR24[11] , 
        \B_DOUT_TEMPR24[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2199 (.A(OR4_2830_Y), .B(OR4_271_Y), .C(OR4_1751_Y), .D(
        OR4_274_Y), .Y(OR4_2199_Y));
    OR4 OR4_484 (.A(\B_DOUT_TEMPR56[38] ), .B(\B_DOUT_TEMPR57[38] ), 
        .C(\B_DOUT_TEMPR58[38] ), .D(\B_DOUT_TEMPR59[38] ), .Y(
        OR4_484_Y));
    OR4 OR4_847 (.A(\A_DOUT_TEMPR79[12] ), .B(\A_DOUT_TEMPR80[12] ), 
        .C(\A_DOUT_TEMPR81[12] ), .D(\A_DOUT_TEMPR82[12] ), .Y(
        OR4_847_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%74%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R74C4 (
        .A_DOUT({nc240, nc241, nc242, nc243, nc244, nc245, nc246, 
        nc247, nc248, nc249, nc250, nc251, nc252, nc253, nc254, 
        \A_DOUT_TEMPR74[24] , \A_DOUT_TEMPR74[23] , 
        \A_DOUT_TEMPR74[22] , \A_DOUT_TEMPR74[21] , 
        \A_DOUT_TEMPR74[20] }), .B_DOUT({nc255, nc256, nc257, nc258, 
        nc259, nc260, nc261, nc262, nc263, nc264, nc265, nc266, nc267, 
        nc268, nc269, \B_DOUT_TEMPR74[24] , \B_DOUT_TEMPR74[23] , 
        \B_DOUT_TEMPR74[22] , \B_DOUT_TEMPR74[21] , 
        \B_DOUT_TEMPR74[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[74][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_616 (.A(OR4_1270_Y), .B(OR4_2150_Y), .C(OR4_1809_Y), .D(
        OR4_266_Y), .Y(OR4_616_Y));
    OR4 OR4_993 (.A(\A_DOUT_TEMPR115[12] ), .B(\A_DOUT_TEMPR116[12] ), 
        .C(\A_DOUT_TEMPR117[12] ), .D(\A_DOUT_TEMPR118[12] ), .Y(
        OR4_993_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[0]  (.A(CFG3_17_Y), .B(
        CFG3_14_Y), .Y(\BLKX2[0] ));
    OR2 OR2_40 (.A(\A_DOUT_TEMPR72[35] ), .B(\A_DOUT_TEMPR73[35] ), .Y(
        OR2_40_Y));
    OR4 OR4_1308 (.A(\B_DOUT_TEMPR48[19] ), .B(\B_DOUT_TEMPR49[19] ), 
        .C(\B_DOUT_TEMPR50[19] ), .D(\B_DOUT_TEMPR51[19] ), .Y(
        OR4_1308_Y));
    OR4 OR4_1666 (.A(OR4_2753_Y), .B(OR4_1132_Y), .C(OR2_17_Y), .D(
        \A_DOUT_TEMPR74[0] ), .Y(OR4_1666_Y));
    OR4 OR4_2030 (.A(\B_DOUT_TEMPR20[23] ), .B(\B_DOUT_TEMPR21[23] ), 
        .C(\B_DOUT_TEMPR22[23] ), .D(\B_DOUT_TEMPR23[23] ), .Y(
        OR4_2030_Y));
    OR4 OR4_2768 (.A(\A_DOUT_TEMPR56[1] ), .B(\A_DOUT_TEMPR57[1] ), .C(
        \A_DOUT_TEMPR58[1] ), .D(\A_DOUT_TEMPR59[1] ), .Y(OR4_2768_Y));
    OR4 \OR4_B_DOUT[36]  (.A(OR4_1103_Y), .B(OR4_3034_Y), .C(OR4_666_Y)
        , .D(OR4_2037_Y), .Y(B_DOUT[36]));
    OR4 OR4_421 (.A(OR4_264_Y), .B(OR4_821_Y), .C(OR4_1507_Y), .D(
        OR4_1800_Y), .Y(OR4_421_Y));
    OR4 OR4_1160 (.A(\A_DOUT_TEMPR52[30] ), .B(\A_DOUT_TEMPR53[30] ), 
        .C(\A_DOUT_TEMPR54[30] ), .D(\A_DOUT_TEMPR55[30] ), .Y(
        OR4_1160_Y));
    OR4 OR4_3010 (.A(\A_DOUT_TEMPR48[22] ), .B(\A_DOUT_TEMPR49[22] ), 
        .C(\A_DOUT_TEMPR50[22] ), .D(\A_DOUT_TEMPR51[22] ), .Y(
        OR4_3010_Y));
    OR4 OR4_2122 (.A(\A_DOUT_TEMPR20[35] ), .B(\A_DOUT_TEMPR21[35] ), 
        .C(\A_DOUT_TEMPR22[35] ), .D(\A_DOUT_TEMPR23[35] ), .Y(
        OR4_2122_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%23%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R23C7 (
        .A_DOUT({nc270, nc271, nc272, nc273, nc274, nc275, nc276, 
        nc277, nc278, nc279, nc280, nc281, nc282, nc283, nc284, 
        \A_DOUT_TEMPR23[39] , \A_DOUT_TEMPR23[38] , 
        \A_DOUT_TEMPR23[37] , \A_DOUT_TEMPR23[36] , 
        \A_DOUT_TEMPR23[35] }), .B_DOUT({nc285, nc286, nc287, nc288, 
        nc289, nc290, nc291, nc292, nc293, nc294, nc295, nc296, nc297, 
        nc298, nc299, \B_DOUT_TEMPR23[39] , \B_DOUT_TEMPR23[38] , 
        \B_DOUT_TEMPR23[37] , \B_DOUT_TEMPR23[36] , 
        \B_DOUT_TEMPR23[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2117 (.A(OR4_1876_Y), .B(OR4_1674_Y), .C(OR2_40_Y), .D(
        \A_DOUT_TEMPR74[35] ), .Y(OR4_2117_Y));
    OR4 OR4_539 (.A(\A_DOUT_TEMPR48[10] ), .B(\A_DOUT_TEMPR49[10] ), 
        .C(\A_DOUT_TEMPR50[10] ), .D(\A_DOUT_TEMPR51[10] ), .Y(
        OR4_539_Y));
    OR4 OR4_1030 (.A(\A_DOUT_TEMPR28[7] ), .B(\A_DOUT_TEMPR29[7] ), .C(
        \A_DOUT_TEMPR30[7] ), .D(\A_DOUT_TEMPR31[7] ), .Y(OR4_1030_Y));
    OR4 OR4_2614 (.A(\B_DOUT_TEMPR64[29] ), .B(\B_DOUT_TEMPR65[29] ), 
        .C(\B_DOUT_TEMPR66[29] ), .D(\B_DOUT_TEMPR67[29] ), .Y(
        OR4_2614_Y));
    OR4 OR4_456 (.A(\A_DOUT_TEMPR52[7] ), .B(\A_DOUT_TEMPR53[7] ), .C(
        \A_DOUT_TEMPR54[7] ), .D(\A_DOUT_TEMPR55[7] ), .Y(OR4_456_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%11%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R11C5 (
        .A_DOUT({nc300, nc301, nc302, nc303, nc304, nc305, nc306, 
        nc307, nc308, nc309, nc310, nc311, nc312, nc313, nc314, 
        \A_DOUT_TEMPR11[29] , \A_DOUT_TEMPR11[28] , 
        \A_DOUT_TEMPR11[27] , \A_DOUT_TEMPR11[26] , 
        \A_DOUT_TEMPR11[25] }), .B_DOUT({nc315, nc316, nc317, nc318, 
        nc319, nc320, nc321, nc322, nc323, nc324, nc325, nc326, nc327, 
        nc328, nc329, \B_DOUT_TEMPR11[29] , \B_DOUT_TEMPR11[28] , 
        \B_DOUT_TEMPR11[27] , \B_DOUT_TEMPR11[26] , 
        \B_DOUT_TEMPR11[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2189 (.A(\A_DOUT_TEMPR52[39] ), .B(\A_DOUT_TEMPR53[39] ), 
        .C(\A_DOUT_TEMPR54[39] ), .D(\A_DOUT_TEMPR55[39] ), .Y(
        OR4_2189_Y));
    OR4 OR4_79 (.A(\A_DOUT_TEMPR16[36] ), .B(\A_DOUT_TEMPR17[36] ), .C(
        \A_DOUT_TEMPR18[36] ), .D(\A_DOUT_TEMPR19[36] ), .Y(OR4_79_Y));
    OR4 \OR4_A_DOUT[33]  (.A(OR4_903_Y), .B(OR4_1397_Y), .C(OR4_585_Y), 
        .D(OR4_1433_Y), .Y(A_DOUT[33]));
    OR4 OR4_1345 (.A(\A_DOUT_TEMPR79[18] ), .B(\A_DOUT_TEMPR80[18] ), 
        .C(\A_DOUT_TEMPR81[18] ), .D(\A_DOUT_TEMPR82[18] ), .Y(
        OR4_1345_Y));
    OR4 OR4_469 (.A(\A_DOUT_TEMPR0[16] ), .B(\A_DOUT_TEMPR1[16] ), .C(
        \A_DOUT_TEMPR2[16] ), .D(\A_DOUT_TEMPR3[16] ), .Y(OR4_469_Y));
    OR4 \OR4_B_DOUT[10]  (.A(OR4_2025_Y), .B(OR4_1445_Y), .C(
        OR4_1186_Y), .D(OR4_2682_Y), .Y(B_DOUT[10]));
    OR4 OR4_114 (.A(OR4_410_Y), .B(OR4_816_Y), .C(OR4_12_Y), .D(
        OR4_1969_Y), .Y(OR4_114_Y));
    OR4 OR4_314 (.A(OR4_2722_Y), .B(OR4_3018_Y), .C(OR4_2645_Y), .D(
        OR4_3036_Y), .Y(OR4_314_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%66%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R66C3 (
        .A_DOUT({nc330, nc331, nc332, nc333, nc334, nc335, nc336, 
        nc337, nc338, nc339, nc340, nc341, nc342, nc343, nc344, 
        \A_DOUT_TEMPR66[19] , \A_DOUT_TEMPR66[18] , 
        \A_DOUT_TEMPR66[17] , \A_DOUT_TEMPR66[16] , 
        \A_DOUT_TEMPR66[15] }), .B_DOUT({nc345, nc346, nc347, nc348, 
        nc349, nc350, nc351, nc352, nc353, nc354, nc355, nc356, nc357, 
        nc358, nc359, \B_DOUT_TEMPR66[19] , \B_DOUT_TEMPR66[18] , 
        \B_DOUT_TEMPR66[17] , \B_DOUT_TEMPR66[16] , 
        \B_DOUT_TEMPR66[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[66][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%4%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R4C3 (
        .A_DOUT({nc360, nc361, nc362, nc363, nc364, nc365, nc366, 
        nc367, nc368, nc369, nc370, nc371, nc372, nc373, nc374, 
        \A_DOUT_TEMPR4[19] , \A_DOUT_TEMPR4[18] , \A_DOUT_TEMPR4[17] , 
        \A_DOUT_TEMPR4[16] , \A_DOUT_TEMPR4[15] }), .B_DOUT({nc375, 
        nc376, nc377, nc378, nc379, nc380, nc381, nc382, nc383, nc384, 
        nc385, nc386, nc387, nc388, nc389, \B_DOUT_TEMPR4[19] , 
        \B_DOUT_TEMPR4[18] , \B_DOUT_TEMPR4[17] , \B_DOUT_TEMPR4[16] , 
        \B_DOUT_TEMPR4[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1027 (.A(\B_DOUT_TEMPR44[10] ), .B(\B_DOUT_TEMPR45[10] ), 
        .C(\B_DOUT_TEMPR46[10] ), .D(\B_DOUT_TEMPR47[10] ), .Y(
        OR4_1027_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%30%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R30C0 (
        .A_DOUT({nc390, nc391, nc392, nc393, nc394, nc395, nc396, 
        nc397, nc398, nc399, nc400, nc401, nc402, nc403, nc404, 
        \A_DOUT_TEMPR30[4] , \A_DOUT_TEMPR30[3] , \A_DOUT_TEMPR30[2] , 
        \A_DOUT_TEMPR30[1] , \A_DOUT_TEMPR30[0] }), .B_DOUT({nc405, 
        nc406, nc407, nc408, nc409, nc410, nc411, nc412, nc413, nc414, 
        nc415, nc416, nc417, nc418, nc419, \B_DOUT_TEMPR30[4] , 
        \B_DOUT_TEMPR30[3] , \B_DOUT_TEMPR30[2] , \B_DOUT_TEMPR30[1] , 
        \B_DOUT_TEMPR30[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2947 (.A(\B_DOUT_TEMPR103[4] ), .B(\B_DOUT_TEMPR104[4] ), 
        .C(\B_DOUT_TEMPR105[4] ), .D(\B_DOUT_TEMPR106[4] ), .Y(
        OR4_2947_Y));
    OR4 OR4_1329 (.A(\A_DOUT_TEMPR91[4] ), .B(\A_DOUT_TEMPR92[4] ), .C(
        \A_DOUT_TEMPR93[4] ), .D(\A_DOUT_TEMPR94[4] ), .Y(OR4_1329_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%35%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R35C4 (
        .A_DOUT({nc420, nc421, nc422, nc423, nc424, nc425, nc426, 
        nc427, nc428, nc429, nc430, nc431, nc432, nc433, nc434, 
        \A_DOUT_TEMPR35[24] , \A_DOUT_TEMPR35[23] , 
        \A_DOUT_TEMPR35[22] , \A_DOUT_TEMPR35[21] , 
        \A_DOUT_TEMPR35[20] }), .B_DOUT({nc435, nc436, nc437, nc438, 
        nc439, nc440, nc441, nc442, nc443, nc444, nc445, nc446, nc447, 
        nc448, nc449, \B_DOUT_TEMPR35[24] , \B_DOUT_TEMPR35[23] , 
        \B_DOUT_TEMPR35[22] , \B_DOUT_TEMPR35[21] , 
        \B_DOUT_TEMPR35[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[35][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1227 (.A(\A_DOUT_TEMPR0[35] ), .B(\A_DOUT_TEMPR1[35] ), .C(
        \A_DOUT_TEMPR2[35] ), .D(\A_DOUT_TEMPR3[35] ), .Y(OR4_1227_Y));
    OR4 OR4_270 (.A(\A_DOUT_TEMPR83[10] ), .B(\A_DOUT_TEMPR84[10] ), 
        .C(\A_DOUT_TEMPR85[10] ), .D(\A_DOUT_TEMPR86[10] ), .Y(
        OR4_270_Y));
    OR4 OR4_670 (.A(\A_DOUT_TEMPR40[1] ), .B(\A_DOUT_TEMPR41[1] ), .C(
        \A_DOUT_TEMPR42[1] ), .D(\A_DOUT_TEMPR43[1] ), .Y(OR4_670_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%58%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R58C6 (
        .A_DOUT({nc450, nc451, nc452, nc453, nc454, nc455, nc456, 
        nc457, nc458, nc459, nc460, nc461, nc462, nc463, nc464, 
        \A_DOUT_TEMPR58[34] , \A_DOUT_TEMPR58[33] , 
        \A_DOUT_TEMPR58[32] , \A_DOUT_TEMPR58[31] , 
        \A_DOUT_TEMPR58[30] }), .B_DOUT({nc465, nc466, nc467, nc468, 
        nc469, nc470, nc471, nc472, nc473, nc474, nc475, nc476, nc477, 
        nc478, nc479, \B_DOUT_TEMPR58[34] , \B_DOUT_TEMPR58[33] , 
        \B_DOUT_TEMPR58[32] , \B_DOUT_TEMPR58[31] , 
        \B_DOUT_TEMPR58[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[58][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2436 (.A(\A_DOUT_TEMPR48[32] ), .B(\A_DOUT_TEMPR49[32] ), 
        .C(\A_DOUT_TEMPR50[32] ), .D(\A_DOUT_TEMPR51[32] ), .Y(
        OR4_2436_Y));
    OR4 OR4_1920 (.A(OR4_2146_Y), .B(OR4_789_Y), .C(OR4_228_Y), .D(
        OR4_1548_Y), .Y(OR4_1920_Y));
    OR4 OR4_1405 (.A(\B_DOUT_TEMPR68[7] ), .B(\B_DOUT_TEMPR69[7] ), .C(
        \B_DOUT_TEMPR70[7] ), .D(\B_DOUT_TEMPR71[7] ), .Y(OR4_1405_Y));
    OR4 OR4_2675 (.A(\B_DOUT_TEMPR40[30] ), .B(\B_DOUT_TEMPR41[30] ), 
        .C(\B_DOUT_TEMPR42[30] ), .D(\B_DOUT_TEMPR43[30] ), .Y(
        OR4_2675_Y));
    OR4 OR4_1179 (.A(\A_DOUT_TEMPR4[5] ), .B(\A_DOUT_TEMPR5[5] ), .C(
        \A_DOUT_TEMPR6[5] ), .D(\A_DOUT_TEMPR7[5] ), .Y(OR4_1179_Y));
    OR4 OR4_161 (.A(\B_DOUT_TEMPR20[29] ), .B(\B_DOUT_TEMPR21[29] ), 
        .C(\B_DOUT_TEMPR22[29] ), .D(\B_DOUT_TEMPR23[29] ), .Y(
        OR4_161_Y));
    OR4 OR4_1094 (.A(OR4_2107_Y), .B(OR4_1578_Y), .C(OR4_2188_Y), .D(
        OR4_1403_Y), .Y(OR4_1094_Y));
    OR4 OR4_1436 (.A(\B_DOUT_TEMPR115[0] ), .B(\B_DOUT_TEMPR116[0] ), 
        .C(\B_DOUT_TEMPR117[0] ), .D(\B_DOUT_TEMPR118[0] ), .Y(
        OR4_1436_Y));
    OR4 OR4_1289 (.A(OR4_2242_Y), .B(OR4_204_Y), .C(OR4_910_Y), .D(
        OR4_2567_Y), .Y(OR4_1289_Y));
    OR4 OR4_1096 (.A(OR4_1758_Y), .B(OR4_2131_Y), .C(OR4_1732_Y), .D(
        OR4_2784_Y), .Y(OR4_1096_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%115%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R115C5 (
        .A_DOUT({nc480, nc481, nc482, nc483, nc484, nc485, nc486, 
        nc487, nc488, nc489, nc490, nc491, nc492, nc493, nc494, 
        \A_DOUT_TEMPR115[29] , \A_DOUT_TEMPR115[28] , 
        \A_DOUT_TEMPR115[27] , \A_DOUT_TEMPR115[26] , 
        \A_DOUT_TEMPR115[25] }), .B_DOUT({nc495, nc496, nc497, nc498, 
        nc499, nc500, nc501, nc502, nc503, nc504, nc505, nc506, nc507, 
        nc508, nc509, \B_DOUT_TEMPR115[29] , \B_DOUT_TEMPR115[28] , 
        \B_DOUT_TEMPR115[27] , \B_DOUT_TEMPR115[26] , 
        \B_DOUT_TEMPR115[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[115][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_884 (.A(\B_DOUT_TEMPR4[6] ), .B(\B_DOUT_TEMPR5[6] ), .C(
        \B_DOUT_TEMPR6[6] ), .D(\B_DOUT_TEMPR7[6] ), .Y(OR4_884_Y));
    OR4 OR4_2840 (.A(\B_DOUT_TEMPR16[36] ), .B(\B_DOUT_TEMPR17[36] ), 
        .C(\B_DOUT_TEMPR18[36] ), .D(\B_DOUT_TEMPR19[36] ), .Y(
        OR4_2840_Y));
    OR4 OR4_441 (.A(\B_DOUT_TEMPR48[26] ), .B(\B_DOUT_TEMPR49[26] ), 
        .C(\B_DOUT_TEMPR50[26] ), .D(\B_DOUT_TEMPR51[26] ), .Y(
        OR4_441_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%23%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R23C0 (
        .A_DOUT({nc510, nc511, nc512, nc513, nc514, nc515, nc516, 
        nc517, nc518, nc519, nc520, nc521, nc522, nc523, nc524, 
        \A_DOUT_TEMPR23[4] , \A_DOUT_TEMPR23[3] , \A_DOUT_TEMPR23[2] , 
        \A_DOUT_TEMPR23[1] , \A_DOUT_TEMPR23[0] }), .B_DOUT({nc525, 
        nc526, nc527, nc528, nc529, nc530, nc531, nc532, nc533, nc534, 
        nc535, nc536, nc537, nc538, nc539, \B_DOUT_TEMPR23[4] , 
        \B_DOUT_TEMPR23[3] , \B_DOUT_TEMPR23[2] , \B_DOUT_TEMPR23[1] , 
        \B_DOUT_TEMPR23[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[25]  (.A(OR4_2628_Y), .B(OR4_2491_Y), .C(
        OR4_1648_Y), .D(OR4_2266_Y), .Y(A_DOUT[25]));
    OR4 OR4_2892 (.A(\B_DOUT_TEMPR115[24] ), .B(\B_DOUT_TEMPR116[24] ), 
        .C(\B_DOUT_TEMPR117[24] ), .D(\B_DOUT_TEMPR118[24] ), .Y(
        OR4_2892_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_6 (.A(B_ADDR[16]), .B(B_ADDR[15]), .C(
        B_ADDR[14]), .Y(CFG3_6_Y));
    OR4 OR4_582 (.A(\B_DOUT_TEMPR115[14] ), .B(\B_DOUT_TEMPR116[14] ), 
        .C(\B_DOUT_TEMPR117[14] ), .D(\B_DOUT_TEMPR118[14] ), .Y(
        OR4_582_Y));
    OR4 OR4_2735 (.A(OR4_1551_Y), .B(OR4_78_Y), .C(OR4_930_Y), .D(
        OR4_2986_Y), .Y(OR4_2735_Y));
    OR4 OR4_1655 (.A(\A_DOUT_TEMPR68[25] ), .B(\A_DOUT_TEMPR69[25] ), 
        .C(\A_DOUT_TEMPR70[25] ), .D(\A_DOUT_TEMPR71[25] ), .Y(
        OR4_1655_Y));
    OR4 OR4_1722 (.A(\B_DOUT_TEMPR64[10] ), .B(\B_DOUT_TEMPR65[10] ), 
        .C(\B_DOUT_TEMPR66[10] ), .D(\B_DOUT_TEMPR67[10] ), .Y(
        OR4_1722_Y));
    OR4 OR4_3 (.A(\A_DOUT_TEMPR87[4] ), .B(\A_DOUT_TEMPR88[4] ), .C(
        \A_DOUT_TEMPR89[4] ), .D(\A_DOUT_TEMPR90[4] ), .Y(OR4_3_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%1%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R1C5 (
        .A_DOUT({nc540, nc541, nc542, nc543, nc544, nc545, nc546, 
        nc547, nc548, nc549, nc550, nc551, nc552, nc553, nc554, 
        \A_DOUT_TEMPR1[29] , \A_DOUT_TEMPR1[28] , \A_DOUT_TEMPR1[27] , 
        \A_DOUT_TEMPR1[26] , \A_DOUT_TEMPR1[25] }), .B_DOUT({nc555, 
        nc556, nc557, nc558, nc559, nc560, nc561, nc562, nc563, nc564, 
        nc565, nc566, nc567, nc568, nc569, \B_DOUT_TEMPR1[29] , 
        \B_DOUT_TEMPR1[28] , \B_DOUT_TEMPR1[27] , \B_DOUT_TEMPR1[26] , 
        \B_DOUT_TEMPR1[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1735 (.A(\A_DOUT_TEMPR8[19] ), .B(\A_DOUT_TEMPR9[19] ), .C(
        \A_DOUT_TEMPR10[19] ), .D(\A_DOUT_TEMPR11[19] ), .Y(OR4_1735_Y)
        );
    OR4 OR4_2844 (.A(\A_DOUT_TEMPR111[18] ), .B(\A_DOUT_TEMPR112[18] ), 
        .C(\A_DOUT_TEMPR113[18] ), .D(\A_DOUT_TEMPR114[18] ), .Y(
        OR4_2844_Y));
    OR4 OR4_2677 (.A(OR4_2157_Y), .B(OR4_456_Y), .C(OR4_93_Y), .D(
        OR4_1177_Y), .Y(OR4_2677_Y));
    OR4 OR4_1393 (.A(\B_DOUT_TEMPR75[27] ), .B(\B_DOUT_TEMPR76[27] ), 
        .C(\B_DOUT_TEMPR77[27] ), .D(\B_DOUT_TEMPR78[27] ), .Y(
        OR4_1393_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[19]  (.A(CFG3_23_Y), .B(
        CFG3_3_Y), .Y(\BLKX2[19] ));
    OR4 OR4_1963 (.A(\B_DOUT_TEMPR20[31] ), .B(\B_DOUT_TEMPR21[31] ), 
        .C(\B_DOUT_TEMPR22[31] ), .D(\B_DOUT_TEMPR23[31] ), .Y(
        OR4_1963_Y));
    OR4 OR4_1706 (.A(\A_DOUT_TEMPR91[37] ), .B(\A_DOUT_TEMPR92[37] ), 
        .C(\A_DOUT_TEMPR93[37] ), .D(\A_DOUT_TEMPR94[37] ), .Y(
        OR4_1706_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%81%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R81C2 (
        .A_DOUT({nc570, nc571, nc572, nc573, nc574, nc575, nc576, 
        nc577, nc578, nc579, nc580, nc581, nc582, nc583, nc584, 
        \A_DOUT_TEMPR81[14] , \A_DOUT_TEMPR81[13] , 
        \A_DOUT_TEMPR81[12] , \A_DOUT_TEMPR81[11] , 
        \A_DOUT_TEMPR81[10] }), .B_DOUT({nc585, nc586, nc587, nc588, 
        nc589, nc590, nc591, nc592, nc593, nc594, nc595, nc596, nc597, 
        nc598, nc599, \B_DOUT_TEMPR81[14] , \B_DOUT_TEMPR81[13] , 
        \B_DOUT_TEMPR81[12] , \B_DOUT_TEMPR81[11] , 
        \B_DOUT_TEMPR81[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[81][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_45 (.A(\A_DOUT_TEMPR72[12] ), .B(\A_DOUT_TEMPR73[12] ), .Y(
        OR2_45_Y));
    OR4 OR4_265 (.A(OR4_3030_Y), .B(OR4_2849_Y), .C(OR4_2801_Y), .D(
        OR4_97_Y), .Y(OR4_265_Y));
    OR4 OR4_200 (.A(\A_DOUT_TEMPR8[28] ), .B(\A_DOUT_TEMPR9[28] ), .C(
        \A_DOUT_TEMPR10[28] ), .D(\A_DOUT_TEMPR11[28] ), .Y(OR4_200_Y));
    OR2 OR2_33 (.A(\B_DOUT_TEMPR72[28] ), .B(\B_DOUT_TEMPR73[28] ), .Y(
        OR2_33_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%27%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R27C7 (
        .A_DOUT({nc600, nc601, nc602, nc603, nc604, nc605, nc606, 
        nc607, nc608, nc609, nc610, nc611, nc612, nc613, nc614, 
        \A_DOUT_TEMPR27[39] , \A_DOUT_TEMPR27[38] , 
        \A_DOUT_TEMPR27[37] , \A_DOUT_TEMPR27[36] , 
        \A_DOUT_TEMPR27[35] }), .B_DOUT({nc615, nc616, nc617, nc618, 
        nc619, nc620, nc621, nc622, nc623, nc624, nc625, nc626, nc627, 
        nc628, nc629, \B_DOUT_TEMPR27[39] , \B_DOUT_TEMPR27[38] , 
        \B_DOUT_TEMPR27[37] , \B_DOUT_TEMPR27[36] , 
        \B_DOUT_TEMPR27[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1513 (.A(OR4_746_Y), .B(OR4_561_Y), .C(OR4_1424_Y), .D(
        OR4_2624_Y), .Y(OR4_1513_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%92%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R92C6 (
        .A_DOUT({nc630, nc631, nc632, nc633, nc634, nc635, nc636, 
        nc637, nc638, nc639, nc640, nc641, nc642, nc643, nc644, 
        \A_DOUT_TEMPR92[34] , \A_DOUT_TEMPR92[33] , 
        \A_DOUT_TEMPR92[32] , \A_DOUT_TEMPR92[31] , 
        \A_DOUT_TEMPR92[30] }), .B_DOUT({nc645, nc646, nc647, nc648, 
        nc649, nc650, nc651, nc652, nc653, nc654, nc655, nc656, nc657, 
        nc658, nc659, \B_DOUT_TEMPR92[34] , \B_DOUT_TEMPR92[33] , 
        \B_DOUT_TEMPR92[32] , \B_DOUT_TEMPR92[31] , 
        \B_DOUT_TEMPR92[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[92][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%54%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R54C3 (
        .A_DOUT({nc660, nc661, nc662, nc663, nc664, nc665, nc666, 
        nc667, nc668, nc669, nc670, nc671, nc672, nc673, nc674, 
        \A_DOUT_TEMPR54[19] , \A_DOUT_TEMPR54[18] , 
        \A_DOUT_TEMPR54[17] , \A_DOUT_TEMPR54[16] , 
        \A_DOUT_TEMPR54[15] }), .B_DOUT({nc675, nc676, nc677, nc678, 
        nc679, nc680, nc681, nc682, nc683, nc684, nc685, nc686, nc687, 
        nc688, nc689, \B_DOUT_TEMPR54[19] , \B_DOUT_TEMPR54[18] , 
        \B_DOUT_TEMPR54[17] , \B_DOUT_TEMPR54[16] , 
        \B_DOUT_TEMPR54[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[54][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_600 (.A(\A_DOUT_TEMPR8[20] ), .B(\A_DOUT_TEMPR9[20] ), .C(
        \A_DOUT_TEMPR10[20] ), .D(\A_DOUT_TEMPR11[20] ), .Y(OR4_600_Y));
    OR4 OR4_2882 (.A(OR4_2586_Y), .B(OR4_2611_Y), .C(OR4_187_Y), .D(
        OR4_2412_Y), .Y(OR4_2882_Y));
    OR4 OR4_2693 (.A(\A_DOUT_TEMPR56[38] ), .B(\A_DOUT_TEMPR57[38] ), 
        .C(\A_DOUT_TEMPR58[38] ), .D(\A_DOUT_TEMPR59[38] ), .Y(
        OR4_2693_Y));
    OR4 OR4_816 (.A(\B_DOUT_TEMPR36[6] ), .B(\B_DOUT_TEMPR37[6] ), .C(
        \B_DOUT_TEMPR38[6] ), .D(\B_DOUT_TEMPR39[6] ), .Y(OR4_816_Y));
    OR4 OR4_2229 (.A(\A_DOUT_TEMPR32[24] ), .B(\A_DOUT_TEMPR33[24] ), 
        .C(\A_DOUT_TEMPR34[24] ), .D(\A_DOUT_TEMPR35[24] ), .Y(
        OR4_2229_Y));
    OR4 OR4_1657 (.A(\B_DOUT_TEMPR28[36] ), .B(\B_DOUT_TEMPR29[36] ), 
        .C(\B_DOUT_TEMPR30[36] ), .D(\B_DOUT_TEMPR31[36] ), .Y(
        OR4_1657_Y));
    OR4 OR4_1113 (.A(\A_DOUT_TEMPR36[1] ), .B(\A_DOUT_TEMPR37[1] ), .C(
        \A_DOUT_TEMPR38[1] ), .D(\A_DOUT_TEMPR39[1] ), .Y(OR4_1113_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%99%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R99C0 (
        .A_DOUT({nc690, nc691, nc692, nc693, nc694, nc695, nc696, 
        nc697, nc698, nc699, nc700, nc701, nc702, nc703, nc704, 
        \A_DOUT_TEMPR99[4] , \A_DOUT_TEMPR99[3] , \A_DOUT_TEMPR99[2] , 
        \A_DOUT_TEMPR99[1] , \A_DOUT_TEMPR99[0] }), .B_DOUT({nc705, 
        nc706, nc707, nc708, nc709, nc710, nc711, nc712, nc713, nc714, 
        nc715, nc716, nc717, nc718, nc719, \B_DOUT_TEMPR99[4] , 
        \B_DOUT_TEMPR99[3] , \B_DOUT_TEMPR99[2] , \B_DOUT_TEMPR99[1] , 
        \B_DOUT_TEMPR99[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[99][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1622 (.A(\A_DOUT_TEMPR4[20] ), .B(\A_DOUT_TEMPR5[20] ), .C(
        \A_DOUT_TEMPR6[20] ), .D(\A_DOUT_TEMPR7[20] ), .Y(OR4_1622_Y));
    OR4 OR4_2610 (.A(\A_DOUT_TEMPR52[10] ), .B(\A_DOUT_TEMPR53[10] ), 
        .C(\A_DOUT_TEMPR54[10] ), .D(\A_DOUT_TEMPR55[10] ), .Y(
        OR4_2610_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%72%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R72C7 (
        .A_DOUT({nc720, nc721, nc722, nc723, nc724, nc725, nc726, 
        nc727, nc728, nc729, nc730, nc731, nc732, nc733, nc734, 
        \A_DOUT_TEMPR72[39] , \A_DOUT_TEMPR72[38] , 
        \A_DOUT_TEMPR72[37] , \A_DOUT_TEMPR72[36] , 
        \A_DOUT_TEMPR72[35] }), .B_DOUT({nc735, nc736, nc737, nc738, 
        nc739, nc740, nc741, nc742, nc743, nc744, nc745, nc746, nc747, 
        nc748, nc749, \B_DOUT_TEMPR72[39] , \B_DOUT_TEMPR72[38] , 
        \B_DOUT_TEMPR72[37] , \B_DOUT_TEMPR72[36] , 
        \B_DOUT_TEMPR72[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[72][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2999 (.A(\A_DOUT_TEMPR24[6] ), .B(\A_DOUT_TEMPR25[6] ), .C(
        \A_DOUT_TEMPR26[6] ), .D(\A_DOUT_TEMPR27[6] ), .Y(OR4_2999_Y));
    OR4 OR4_1361 (.A(\A_DOUT_TEMPR44[4] ), .B(\A_DOUT_TEMPR45[4] ), .C(
        \A_DOUT_TEMPR46[4] ), .D(\A_DOUT_TEMPR47[4] ), .Y(OR4_1361_Y));
    OR4 OR4_666 (.A(OR4_305_Y), .B(OR4_1253_Y), .C(OR4_897_Y), .D(
        OR4_2369_Y), .Y(OR4_666_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%38%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R38C6 (
        .A_DOUT({nc750, nc751, nc752, nc753, nc754, nc755, nc756, 
        nc757, nc758, nc759, nc760, nc761, nc762, nc763, nc764, 
        \A_DOUT_TEMPR38[34] , \A_DOUT_TEMPR38[33] , 
        \A_DOUT_TEMPR38[32] , \A_DOUT_TEMPR38[31] , 
        \A_DOUT_TEMPR38[30] }), .B_DOUT({nc765, nc766, nc767, nc768, 
        nc769, nc770, nc771, nc772, nc773, nc774, nc775, nc776, nc777, 
        nc778, nc779, \B_DOUT_TEMPR38[34] , \B_DOUT_TEMPR38[33] , 
        \B_DOUT_TEMPR38[32] , \B_DOUT_TEMPR38[31] , 
        \B_DOUT_TEMPR38[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[38][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_829 (.A(OR4_1508_Y), .B(OR4_1890_Y), .C(OR4_1486_Y), .D(
        OR4_2505_Y), .Y(OR4_829_Y));
    OR4 OR4_496 (.A(\B_DOUT_TEMPR24[5] ), .B(\B_DOUT_TEMPR25[5] ), .C(
        \B_DOUT_TEMPR26[5] ), .D(\B_DOUT_TEMPR27[5] ), .Y(OR4_496_Y));
    OR4 OR4_310 (.A(\A_DOUT_TEMPR52[32] ), .B(\A_DOUT_TEMPR53[32] ), 
        .C(\A_DOUT_TEMPR54[32] ), .D(\A_DOUT_TEMPR55[32] ), .Y(
        OR4_310_Y));
    OR4 OR4_2018 (.A(\B_DOUT_TEMPR20[15] ), .B(\B_DOUT_TEMPR21[15] ), 
        .C(\B_DOUT_TEMPR22[15] ), .D(\B_DOUT_TEMPR23[15] ), .Y(
        OR4_2018_Y));
    OR4 OR4_1861 (.A(\A_DOUT_TEMPR56[39] ), .B(\A_DOUT_TEMPR57[39] ), 
        .C(\A_DOUT_TEMPR58[39] ), .D(\A_DOUT_TEMPR59[39] ), .Y(
        OR4_1861_Y));
    OR4 OR4_1012 (.A(\A_DOUT_TEMPR8[21] ), .B(\A_DOUT_TEMPR9[21] ), .C(
        \A_DOUT_TEMPR10[21] ), .D(\A_DOUT_TEMPR11[21] ), .Y(OR4_1012_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%118%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R118C7 (
        .A_DOUT({nc780, nc781, nc782, nc783, nc784, nc785, nc786, 
        nc787, nc788, nc789, nc790, nc791, nc792, nc793, nc794, 
        \A_DOUT_TEMPR118[39] , \A_DOUT_TEMPR118[38] , 
        \A_DOUT_TEMPR118[37] , \A_DOUT_TEMPR118[36] , 
        \A_DOUT_TEMPR118[35] }), .B_DOUT({nc795, nc796, nc797, nc798, 
        nc799, nc800, nc801, nc802, nc803, nc804, nc805, nc806, nc807, 
        nc808, nc809, \B_DOUT_TEMPR118[39] , \B_DOUT_TEMPR118[38] , 
        \B_DOUT_TEMPR118[37] , \B_DOUT_TEMPR118[36] , 
        \B_DOUT_TEMPR118[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[118][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[24]  (.A(CFG3_11_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[24] ));
    OR4 OR4_1922 (.A(\A_DOUT_TEMPR36[12] ), .B(\A_DOUT_TEMPR37[12] ), 
        .C(\A_DOUT_TEMPR38[12] ), .D(\A_DOUT_TEMPR39[12] ), .Y(
        OR4_1922_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%95%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R95C6 (
        .A_DOUT({nc810, nc811, nc812, nc813, nc814, nc815, nc816, 
        nc817, nc818, nc819, nc820, nc821, nc822, nc823, nc824, 
        \A_DOUT_TEMPR95[34] , \A_DOUT_TEMPR95[33] , 
        \A_DOUT_TEMPR95[32] , \A_DOUT_TEMPR95[31] , 
        \A_DOUT_TEMPR95[30] }), .B_DOUT({nc825, nc826, nc827, nc828, 
        nc829, nc830, nc831, nc832, nc833, nc834, nc835, nc836, nc837, 
        nc838, nc839, \B_DOUT_TEMPR95[34] , \B_DOUT_TEMPR95[33] , 
        \B_DOUT_TEMPR95[32] , \B_DOUT_TEMPR95[31] , 
        \B_DOUT_TEMPR95[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[95][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_433 (.A(\A_DOUT_TEMPR64[10] ), .B(\A_DOUT_TEMPR65[10] ), 
        .C(\A_DOUT_TEMPR66[10] ), .D(\A_DOUT_TEMPR67[10] ), .Y(
        OR4_433_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%48%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R48C1 (
        .A_DOUT({nc840, nc841, nc842, nc843, nc844, nc845, nc846, 
        nc847, nc848, nc849, nc850, nc851, nc852, nc853, nc854, 
        \A_DOUT_TEMPR48[9] , \A_DOUT_TEMPR48[8] , \A_DOUT_TEMPR48[7] , 
        \A_DOUT_TEMPR48[6] , \A_DOUT_TEMPR48[5] }), .B_DOUT({nc855, 
        nc856, nc857, nc858, nc859, nc860, nc861, nc862, nc863, nc864, 
        nc865, nc866, nc867, nc868, nc869, \B_DOUT_TEMPR48[9] , 
        \B_DOUT_TEMPR48[8] , \B_DOUT_TEMPR48[7] , \B_DOUT_TEMPR48[6] , 
        \B_DOUT_TEMPR48[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[48][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_221 (.A(OR4_1702_Y), .B(OR4_158_Y), .C(OR4_747_Y), .D(
        OR4_566_Y), .Y(OR4_221_Y));
    OR4 OR4_821 (.A(\A_DOUT_TEMPR75[38] ), .B(\A_DOUT_TEMPR76[38] ), 
        .C(\A_DOUT_TEMPR77[38] ), .D(\A_DOUT_TEMPR78[38] ), .Y(
        OR4_821_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%48%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R48C7 (
        .A_DOUT({nc870, nc871, nc872, nc873, nc874, nc875, nc876, 
        nc877, nc878, nc879, nc880, nc881, nc882, nc883, nc884, 
        \A_DOUT_TEMPR48[39] , \A_DOUT_TEMPR48[38] , 
        \A_DOUT_TEMPR48[37] , \A_DOUT_TEMPR48[36] , 
        \A_DOUT_TEMPR48[35] }), .B_DOUT({nc885, nc886, nc887, nc888, 
        nc889, nc890, nc891, nc892, nc893, nc894, nc895, nc896, nc897, 
        nc898, nc899, \B_DOUT_TEMPR48[39] , \B_DOUT_TEMPR48[38] , 
        \B_DOUT_TEMPR48[37] , \B_DOUT_TEMPR48[36] , 
        \B_DOUT_TEMPR48[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[48][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2553 (.A(\B_DOUT_TEMPR28[13] ), .B(\B_DOUT_TEMPR29[13] ), 
        .C(\B_DOUT_TEMPR30[13] ), .D(\B_DOUT_TEMPR31[13] ), .Y(
        OR4_2553_Y));
    OR4 OR4_62 (.A(\A_DOUT_TEMPR79[14] ), .B(\A_DOUT_TEMPR80[14] ), .C(
        \A_DOUT_TEMPR81[14] ), .D(\A_DOUT_TEMPR82[14] ), .Y(OR4_62_Y));
    OR4 OR4_2683 (.A(OR4_1987_Y), .B(OR4_2275_Y), .C(OR4_1927_Y), .D(
        OR4_2294_Y), .Y(OR4_2683_Y));
    OR4 OR4_2794 (.A(\B_DOUT_TEMPR24[23] ), .B(\B_DOUT_TEMPR25[23] ), 
        .C(\B_DOUT_TEMPR26[23] ), .D(\B_DOUT_TEMPR27[23] ), .Y(
        OR4_2794_Y));
    OR4 OR4_2169 (.A(OR4_1277_Y), .B(OR4_592_Y), .C(OR4_2508_Y), .D(
        OR4_731_Y), .Y(OR4_2169_Y));
    OR4 OR4_2989 (.A(\A_DOUT_TEMPR56[9] ), .B(\A_DOUT_TEMPR57[9] ), .C(
        \A_DOUT_TEMPR58[9] ), .D(\A_DOUT_TEMPR59[9] ), .Y(OR4_2989_Y));
    OR4 OR4_2153 (.A(OR4_1691_Y), .B(OR4_1427_Y), .C(OR4_2123_Y), .D(
        OR4_2414_Y), .Y(OR4_2153_Y));
    OR4 OR4_2491 (.A(OR4_733_Y), .B(OR4_1955_Y), .C(OR4_2602_Y), .D(
        OR4_1763_Y), .Y(OR4_2491_Y));
    OR4 OR4_1872 (.A(\B_DOUT_TEMPR103[22] ), .B(\B_DOUT_TEMPR104[22] ), 
        .C(\B_DOUT_TEMPR105[22] ), .D(\B_DOUT_TEMPR106[22] ), .Y(
        OR4_1872_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%82%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R82C3 (
        .A_DOUT({nc900, nc901, nc902, nc903, nc904, nc905, nc906, 
        nc907, nc908, nc909, nc910, nc911, nc912, nc913, nc914, 
        \A_DOUT_TEMPR82[19] , \A_DOUT_TEMPR82[18] , 
        \A_DOUT_TEMPR82[17] , \A_DOUT_TEMPR82[16] , 
        \A_DOUT_TEMPR82[15] }), .B_DOUT({nc915, nc916, nc917, nc918, 
        nc919, nc920, nc921, nc922, nc923, nc924, nc925, nc926, nc927, 
        nc928, nc929, \B_DOUT_TEMPR82[19] , \B_DOUT_TEMPR82[18] , 
        \B_DOUT_TEMPR82[17] , \B_DOUT_TEMPR82[16] , 
        \B_DOUT_TEMPR82[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[82][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2374 (.A(OR4_418_Y), .B(OR4_1836_Y), .C(OR4_1352_Y), .D(
        OR4_1613_Y), .Y(OR4_2374_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%16%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R16C3 (
        .A_DOUT({nc930, nc931, nc932, nc933, nc934, nc935, nc936, 
        nc937, nc938, nc939, nc940, nc941, nc942, nc943, nc944, 
        \A_DOUT_TEMPR16[19] , \A_DOUT_TEMPR16[18] , 
        \A_DOUT_TEMPR16[17] , \A_DOUT_TEMPR16[16] , 
        \A_DOUT_TEMPR16[15] }), .B_DOUT({nc945, nc946, nc947, nc948, 
        nc949, nc950, nc951, nc952, nc953, nc954, nc955, nc956, nc957, 
        nc958, nc959, \B_DOUT_TEMPR16[19] , \B_DOUT_TEMPR16[18] , 
        \B_DOUT_TEMPR16[17] , \B_DOUT_TEMPR16[16] , 
        \B_DOUT_TEMPR16[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2052 (.A(\A_DOUT_TEMPR56[27] ), .B(\A_DOUT_TEMPR57[27] ), 
        .C(\A_DOUT_TEMPR58[27] ), .D(\A_DOUT_TEMPR59[27] ), .Y(
        OR4_2052_Y));
    OR4 OR4_164 (.A(\B_DOUT_TEMPR87[27] ), .B(\B_DOUT_TEMPR88[27] ), 
        .C(\B_DOUT_TEMPR89[27] ), .D(\B_DOUT_TEMPR90[27] ), .Y(
        OR4_164_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%80%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R80C3 (
        .A_DOUT({nc960, nc961, nc962, nc963, nc964, nc965, nc966, 
        nc967, nc968, nc969, nc970, nc971, nc972, nc973, nc974, 
        \A_DOUT_TEMPR80[19] , \A_DOUT_TEMPR80[18] , 
        \A_DOUT_TEMPR80[17] , \A_DOUT_TEMPR80[16] , 
        \A_DOUT_TEMPR80[15] }), .B_DOUT({nc975, nc976, nc977, nc978, 
        nc979, nc980, nc981, nc982, nc983, nc984, nc985, nc986, nc987, 
        nc988, nc989, \B_DOUT_TEMPR80[19] , \B_DOUT_TEMPR80[18] , 
        \B_DOUT_TEMPR80[17] , \B_DOUT_TEMPR80[16] , 
        \B_DOUT_TEMPR80[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[80][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_8 (.A(\A_DOUT_TEMPR52[38] ), .B(\A_DOUT_TEMPR53[38] ), .C(
        \A_DOUT_TEMPR54[38] ), .D(\A_DOUT_TEMPR55[38] ), .Y(OR4_8_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%60%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R60C0 (
        .A_DOUT({nc990, nc991, nc992, nc993, nc994, nc995, nc996, 
        nc997, nc998, nc999, nc1000, nc1001, nc1002, nc1003, nc1004, 
        \A_DOUT_TEMPR60[4] , \A_DOUT_TEMPR60[3] , \A_DOUT_TEMPR60[2] , 
        \A_DOUT_TEMPR60[1] , \A_DOUT_TEMPR60[0] }), .B_DOUT({nc1005, 
        nc1006, nc1007, nc1008, nc1009, nc1010, nc1011, nc1012, nc1013, 
        nc1014, nc1015, nc1016, nc1017, nc1018, nc1019, 
        \B_DOUT_TEMPR60[4] , \B_DOUT_TEMPR60[3] , \B_DOUT_TEMPR60[2] , 
        \B_DOUT_TEMPR60[1] , \B_DOUT_TEMPR60[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[60][0] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[4], 
        B_DIN[3], B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_364 (.A(\A_DOUT_TEMPR48[6] ), .B(\A_DOUT_TEMPR49[6] ), .C(
        \A_DOUT_TEMPR50[6] ), .D(\A_DOUT_TEMPR51[6] ), .Y(OR4_364_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%65%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R65C4 (
        .A_DOUT({nc1020, nc1021, nc1022, nc1023, nc1024, nc1025, 
        nc1026, nc1027, nc1028, nc1029, nc1030, nc1031, nc1032, nc1033, 
        nc1034, \A_DOUT_TEMPR65[24] , \A_DOUT_TEMPR65[23] , 
        \A_DOUT_TEMPR65[22] , \A_DOUT_TEMPR65[21] , 
        \A_DOUT_TEMPR65[20] }), .B_DOUT({nc1035, nc1036, nc1037, 
        nc1038, nc1039, nc1040, nc1041, nc1042, nc1043, nc1044, nc1045, 
        nc1046, nc1047, nc1048, nc1049, \B_DOUT_TEMPR65[24] , 
        \B_DOUT_TEMPR65[23] , \B_DOUT_TEMPR65[22] , 
        \B_DOUT_TEMPR65[21] , \B_DOUT_TEMPR65[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[65][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h2) )  CFG3_12 (.A(B_ADDR[16]), .B(B_ADDR[15]), .C(
        B_ADDR[14]), .Y(CFG3_12_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%34%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R34C3 (
        .A_DOUT({nc1050, nc1051, nc1052, nc1053, nc1054, nc1055, 
        nc1056, nc1057, nc1058, nc1059, nc1060, nc1061, nc1062, nc1063, 
        nc1064, \A_DOUT_TEMPR34[19] , \A_DOUT_TEMPR34[18] , 
        \A_DOUT_TEMPR34[17] , \A_DOUT_TEMPR34[16] , 
        \A_DOUT_TEMPR34[15] }), .B_DOUT({nc1065, nc1066, nc1067, 
        nc1068, nc1069, nc1070, nc1071, nc1072, nc1073, nc1074, nc1075, 
        nc1076, nc1077, nc1078, nc1079, \B_DOUT_TEMPR34[19] , 
        \B_DOUT_TEMPR34[18] , \B_DOUT_TEMPR34[17] , 
        \B_DOUT_TEMPR34[16] , \B_DOUT_TEMPR34[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[34][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2114 (.A(\B_DOUT_TEMPR87[7] ), .B(\B_DOUT_TEMPR88[7] ), .C(
        \B_DOUT_TEMPR89[7] ), .D(\B_DOUT_TEMPR90[7] ), .Y(OR4_2114_Y));
    OR4 OR4_2536 (.A(OR4_404_Y), .B(OR4_1592_Y), .C(OR4_2653_Y), .D(
        OR4_2594_Y), .Y(OR4_2536_Y));
    OR4 OR4_2784 (.A(OR4_551_Y), .B(OR4_2617_Y), .C(OR4_2838_Y), .D(
        OR4_2629_Y), .Y(OR4_2784_Y));
    OR4 OR4_2737 (.A(\B_DOUT_TEMPR79[26] ), .B(\B_DOUT_TEMPR80[26] ), 
        .C(\B_DOUT_TEMPR81[26] ), .D(\B_DOUT_TEMPR82[26] ), .Y(
        OR4_2737_Y));
    OR4 \OR4_A_DOUT[36]  (.A(OR4_2689_Y), .B(OR4_277_Y), .C(OR4_2078_Y)
        , .D(OR4_2093_Y), .Y(A_DOUT[36]));
    OR4 OR4_1354 (.A(\B_DOUT_TEMPR83[6] ), .B(\B_DOUT_TEMPR84[6] ), .C(
        \B_DOUT_TEMPR85[6] ), .D(\B_DOUT_TEMPR86[6] ), .Y(OR4_1354_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%86%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R86C6 (
        .A_DOUT({nc1080, nc1081, nc1082, nc1083, nc1084, nc1085, 
        nc1086, nc1087, nc1088, nc1089, nc1090, nc1091, nc1092, nc1093, 
        nc1094, \A_DOUT_TEMPR86[34] , \A_DOUT_TEMPR86[33] , 
        \A_DOUT_TEMPR86[32] , \A_DOUT_TEMPR86[31] , 
        \A_DOUT_TEMPR86[30] }), .B_DOUT({nc1095, nc1096, nc1097, 
        nc1098, nc1099, nc1100, nc1101, nc1102, nc1103, nc1104, nc1105, 
        nc1106, nc1107, nc1108, nc1109, \B_DOUT_TEMPR86[34] , 
        \B_DOUT_TEMPR86[33] , \B_DOUT_TEMPR86[32] , 
        \B_DOUT_TEMPR86[31] , \B_DOUT_TEMPR86[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[86][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2481 (.A(\A_DOUT_TEMPR91[13] ), .B(\A_DOUT_TEMPR92[13] ), 
        .C(\A_DOUT_TEMPR93[13] ), .D(\A_DOUT_TEMPR94[13] ), .Y(
        OR4_2481_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%9%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R9C5 (
        .A_DOUT({nc1110, nc1111, nc1112, nc1113, nc1114, nc1115, 
        nc1116, nc1117, nc1118, nc1119, nc1120, nc1121, nc1122, nc1123, 
        nc1124, \A_DOUT_TEMPR9[29] , \A_DOUT_TEMPR9[28] , 
        \A_DOUT_TEMPR9[27] , \A_DOUT_TEMPR9[26] , \A_DOUT_TEMPR9[25] })
        , .B_DOUT({nc1125, nc1126, nc1127, nc1128, nc1129, nc1130, 
        nc1131, nc1132, nc1133, nc1134, nc1135, nc1136, nc1137, nc1138, 
        nc1139, \B_DOUT_TEMPR9[29] , \B_DOUT_TEMPR9[28] , 
        \B_DOUT_TEMPR9[27] , \B_DOUT_TEMPR9[26] , \B_DOUT_TEMPR9[25] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[9][5] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[29], A_DIN[28], A_DIN[27], 
        A_DIN[26], A_DIN[25]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1536 (.A(\B_DOUT_TEMPR111[28] ), .B(\B_DOUT_TEMPR112[28] ), 
        .C(\B_DOUT_TEMPR113[28] ), .D(\B_DOUT_TEMPR114[28] ), .Y(
        OR4_1536_Y));
    OR4 OR4_2531 (.A(OR4_774_Y), .B(OR4_1100_Y), .C(OR4_713_Y), .D(
        OR4_1118_Y), .Y(OR4_2531_Y));
    OR4 OR4_1507 (.A(\A_DOUT_TEMPR79[38] ), .B(\A_DOUT_TEMPR80[38] ), 
        .C(\A_DOUT_TEMPR81[38] ), .D(\A_DOUT_TEMPR82[38] ), .Y(
        OR4_1507_Y));
    OR4 OR4_1673 (.A(\A_DOUT_TEMPR95[14] ), .B(\A_DOUT_TEMPR96[14] ), 
        .C(\A_DOUT_TEMPR97[14] ), .D(\A_DOUT_TEMPR98[14] ), .Y(
        OR4_1673_Y));
    OR4 OR4_327 (.A(OR4_2433_Y), .B(OR4_1622_Y), .C(OR4_600_Y), .D(
        OR4_922_Y), .Y(OR4_327_Y));
    OR4 OR4_849 (.A(\B_DOUT_TEMPR87[1] ), .B(\B_DOUT_TEMPR88[1] ), .C(
        \B_DOUT_TEMPR89[1] ), .D(\B_DOUT_TEMPR90[1] ), .Y(OR4_849_Y));
    OR4 OR4_1737 (.A(\B_DOUT_TEMPR111[22] ), .B(\B_DOUT_TEMPR112[22] ), 
        .C(\B_DOUT_TEMPR113[22] ), .D(\B_DOUT_TEMPR114[22] ), .Y(
        OR4_1737_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[26]  (.A(CFG3_22_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[26] ));
    OR4 OR4_2994 (.A(\B_DOUT_TEMPR52[8] ), .B(\B_DOUT_TEMPR53[8] ), .C(
        \B_DOUT_TEMPR54[8] ), .D(\B_DOUT_TEMPR55[8] ), .Y(OR4_2994_Y));
    OR4 OR4_1979 (.A(OR4_2197_Y), .B(OR4_872_Y), .C(OR4_288_Y), .D(
        OR4_1610_Y), .Y(OR4_1979_Y));
    OR4 OR4_250 (.A(OR4_149_Y), .B(OR4_1821_Y), .C(OR4_1229_Y), .D(
        OR4_534_Y), .Y(OR4_250_Y));
    OR4 OR4_1531 (.A(\B_DOUT_TEMPR64[28] ), .B(\B_DOUT_TEMPR65[28] ), 
        .C(\B_DOUT_TEMPR66[28] ), .D(\B_DOUT_TEMPR67[28] ), .Y(
        OR4_1531_Y));
    OR4 OR4_2345 (.A(OR4_2203_Y), .B(OR4_683_Y), .C(OR4_245_Y), .D(
        OR4_1932_Y), .Y(OR4_2345_Y));
    OR4 OR4_828 (.A(OR4_1826_Y), .B(OR4_109_Y), .C(OR4_2817_Y), .D(
        OR4_813_Y), .Y(OR4_828_Y));
    OR4 OR4_241 (.A(\B_DOUT_TEMPR56[17] ), .B(\B_DOUT_TEMPR57[17] ), 
        .C(\B_DOUT_TEMPR58[17] ), .D(\B_DOUT_TEMPR59[17] ), .Y(
        OR4_241_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%41%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R41C1 (
        .A_DOUT({nc1140, nc1141, nc1142, nc1143, nc1144, nc1145, 
        nc1146, nc1147, nc1148, nc1149, nc1150, nc1151, nc1152, nc1153, 
        nc1154, \A_DOUT_TEMPR41[9] , \A_DOUT_TEMPR41[8] , 
        \A_DOUT_TEMPR41[7] , \A_DOUT_TEMPR41[6] , \A_DOUT_TEMPR41[5] })
        , .B_DOUT({nc1155, nc1156, nc1157, nc1158, nc1159, nc1160, 
        nc1161, nc1162, nc1163, nc1164, nc1165, nc1166, nc1167, nc1168, 
        nc1169, \B_DOUT_TEMPR41[9] , \B_DOUT_TEMPR41[8] , 
        \B_DOUT_TEMPR41[7] , \B_DOUT_TEMPR41[6] , \B_DOUT_TEMPR41[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[41][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_621 (.A(\A_DOUT_TEMPR8[33] ), .B(\A_DOUT_TEMPR9[33] ), .C(
        \A_DOUT_TEMPR10[33] ), .D(\A_DOUT_TEMPR11[33] ), .Y(OR4_621_Y));
    OR4 OR4_841 (.A(\A_DOUT_TEMPR56[19] ), .B(\A_DOUT_TEMPR57[19] ), 
        .C(\A_DOUT_TEMPR58[19] ), .D(\A_DOUT_TEMPR59[19] ), .Y(
        OR4_841_Y));
    OR4 OR4_1429 (.A(\A_DOUT_TEMPR64[23] ), .B(\A_DOUT_TEMPR65[23] ), 
        .C(\A_DOUT_TEMPR66[23] ), .D(\A_DOUT_TEMPR67[23] ), .Y(
        OR4_1429_Y));
    OR4 OR4_650 (.A(OR4_1248_Y), .B(OR4_559_Y), .C(OR2_62_Y), .D(
        \B_DOUT_TEMPR74[2] ), .Y(OR4_650_Y));
    OR2 OR2_49 (.A(\A_DOUT_TEMPR72[6] ), .B(\A_DOUT_TEMPR73[6] ), .Y(
        OR2_49_Y));
    OR4 OR4_1543 (.A(OR4_15_Y), .B(OR4_386_Y), .C(OR4_1147_Y), .D(
        OR4_1951_Y), .Y(OR4_1543_Y));
    OR4 OR4_2996 (.A(\B_DOUT_TEMPR20[17] ), .B(\B_DOUT_TEMPR21[17] ), 
        .C(\B_DOUT_TEMPR22[17] ), .D(\B_DOUT_TEMPR23[17] ), .Y(
        OR4_2996_Y));
    OR4 OR4_214 (.A(\B_DOUT_TEMPR12[39] ), .B(\B_DOUT_TEMPR13[39] ), 
        .C(\B_DOUT_TEMPR14[39] ), .D(\B_DOUT_TEMPR15[39] ), .Y(
        OR4_214_Y));
    OR4 OR4_64 (.A(\A_DOUT_TEMPR8[35] ), .B(\A_DOUT_TEMPR9[35] ), .C(
        \A_DOUT_TEMPR10[35] ), .D(\A_DOUT_TEMPR11[35] ), .Y(OR4_64_Y));
    OR4 OR4_2815 (.A(\A_DOUT_TEMPR24[17] ), .B(\A_DOUT_TEMPR25[17] ), 
        .C(\A_DOUT_TEMPR26[17] ), .D(\A_DOUT_TEMPR27[17] ), .Y(
        OR4_2815_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[10]  (.A(CFG3_22_Y), .B(
        CFG3_15_Y), .Y(\BLKY2[10] ));
    OR4 OR4_1143 (.A(\A_DOUT_TEMPR4[27] ), .B(\A_DOUT_TEMPR5[27] ), .C(
        \A_DOUT_TEMPR6[27] ), .D(\A_DOUT_TEMPR7[27] ), .Y(OR4_1143_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%106%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R106C2 (
        .A_DOUT({nc1170, nc1171, nc1172, nc1173, nc1174, nc1175, 
        nc1176, nc1177, nc1178, nc1179, nc1180, nc1181, nc1182, nc1183, 
        nc1184, \A_DOUT_TEMPR106[14] , \A_DOUT_TEMPR106[13] , 
        \A_DOUT_TEMPR106[12] , \A_DOUT_TEMPR106[11] , 
        \A_DOUT_TEMPR106[10] }), .B_DOUT({nc1185, nc1186, nc1187, 
        nc1188, nc1189, nc1190, nc1191, nc1192, nc1193, nc1194, nc1195, 
        nc1196, nc1197, nc1198, nc1199, \B_DOUT_TEMPR106[14] , 
        \B_DOUT_TEMPR106[13] , \B_DOUT_TEMPR106[12] , 
        \B_DOUT_TEMPR106[11] , \B_DOUT_TEMPR106[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[106][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_42 (.A(\B_DOUT_TEMPR64[35] ), .B(\B_DOUT_TEMPR65[35] ), .C(
        \B_DOUT_TEMPR66[35] ), .D(\B_DOUT_TEMPR67[35] ), .Y(OR4_42_Y));
    OR4 OR4_710 (.A(\A_DOUT_TEMPR68[39] ), .B(\A_DOUT_TEMPR69[39] ), 
        .C(\A_DOUT_TEMPR70[39] ), .D(\A_DOUT_TEMPR71[39] ), .Y(
        OR4_710_Y));
    OR4 OR4_1042 (.A(\A_DOUT_TEMPR0[15] ), .B(\A_DOUT_TEMPR1[15] ), .C(
        \A_DOUT_TEMPR2[15] ), .D(\A_DOUT_TEMPR3[15] ), .Y(OR4_1042_Y));
    OR4 OR4_1774 (.A(\A_DOUT_TEMPR56[29] ), .B(\A_DOUT_TEMPR57[29] ), 
        .C(\A_DOUT_TEMPR58[29] ), .D(\A_DOUT_TEMPR59[29] ), .Y(
        OR4_1774_Y));
    OR4 OR4_424 (.A(\B_DOUT_TEMPR48[35] ), .B(\B_DOUT_TEMPR49[35] ), 
        .C(\B_DOUT_TEMPR50[35] ), .D(\B_DOUT_TEMPR51[35] ), .Y(
        OR4_424_Y));
    OR4 OR4_2984 (.A(\A_DOUT_TEMPR52[28] ), .B(\A_DOUT_TEMPR53[28] ), 
        .C(\A_DOUT_TEMPR54[28] ), .D(\A_DOUT_TEMPR55[28] ), .Y(
        OR4_2984_Y));
    OR4 OR4_1981 (.A(\A_DOUT_TEMPR56[12] ), .B(\A_DOUT_TEMPR57[12] ), 
        .C(\A_DOUT_TEMPR58[12] ), .D(\A_DOUT_TEMPR59[12] ), .Y(
        OR4_1981_Y));
    OR4 OR4_1471 (.A(\A_DOUT_TEMPR91[14] ), .B(\A_DOUT_TEMPR92[14] ), 
        .C(\A_DOUT_TEMPR93[14] ), .D(\A_DOUT_TEMPR94[14] ), .Y(
        OR4_1471_Y));
    OR4 OR4_1320 (.A(\B_DOUT_TEMPR79[11] ), .B(\B_DOUT_TEMPR80[11] ), 
        .C(\B_DOUT_TEMPR81[11] ), .D(\B_DOUT_TEMPR82[11] ), .Y(
        OR4_1320_Y));
    OR4 OR4_1427 (.A(\B_DOUT_TEMPR36[39] ), .B(\B_DOUT_TEMPR37[39] ), 
        .C(\B_DOUT_TEMPR38[39] ), .D(\B_DOUT_TEMPR39[39] ), .Y(
        OR4_1427_Y));
    OR4 OR4_2986 (.A(\B_DOUT_TEMPR12[17] ), .B(\B_DOUT_TEMPR13[17] ), 
        .C(\B_DOUT_TEMPR14[17] ), .D(\B_DOUT_TEMPR15[17] ), .Y(
        OR4_2986_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENB[10]  (.A(B_WBYTE_EN[5]), .B(
        B_WEN), .Y(\WBYTEENB[10] ));
    OR4 OR4_866 (.A(OR4_42_Y), .B(OR4_2906_Y), .C(OR2_73_Y), .D(
        \B_DOUT_TEMPR74[35] ), .Y(OR4_866_Y));
    OR4 OR4_2862 (.A(\A_DOUT_TEMPR103[35] ), .B(\A_DOUT_TEMPR104[35] ), 
        .C(\A_DOUT_TEMPR105[35] ), .D(\A_DOUT_TEMPR106[35] ), .Y(
        OR4_2862_Y));
    OR4 OR4_2470 (.A(\B_DOUT_TEMPR40[10] ), .B(\B_DOUT_TEMPR41[10] ), 
        .C(\B_DOUT_TEMPR42[10] ), .D(\B_DOUT_TEMPR43[10] ), .Y(
        OR4_2470_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%110%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R110C3 (
        .A_DOUT({nc1200, nc1201, nc1202, nc1203, nc1204, nc1205, 
        nc1206, nc1207, nc1208, nc1209, nc1210, nc1211, nc1212, nc1213, 
        nc1214, \A_DOUT_TEMPR110[19] , \A_DOUT_TEMPR110[18] , 
        \A_DOUT_TEMPR110[17] , \A_DOUT_TEMPR110[16] , 
        \A_DOUT_TEMPR110[15] }), .B_DOUT({nc1215, nc1216, nc1217, 
        nc1218, nc1219, nc1220, nc1221, nc1222, nc1223, nc1224, nc1225, 
        nc1226, nc1227, nc1228, nc1229, \B_DOUT_TEMPR110[19] , 
        \B_DOUT_TEMPR110[18] , \B_DOUT_TEMPR110[17] , 
        \B_DOUT_TEMPR110[16] , \B_DOUT_TEMPR110[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[110][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_3034 (.A(OR4_2482_Y), .B(OR4_756_Y), .C(OR4_1449_Y), .D(
        OR4_1744_Y), .Y(OR4_3034_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%68%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R68C6 (
        .A_DOUT({nc1230, nc1231, nc1232, nc1233, nc1234, nc1235, 
        nc1236, nc1237, nc1238, nc1239, nc1240, nc1241, nc1242, nc1243, 
        nc1244, \A_DOUT_TEMPR68[34] , \A_DOUT_TEMPR68[33] , 
        \A_DOUT_TEMPR68[32] , \A_DOUT_TEMPR68[31] , 
        \A_DOUT_TEMPR68[30] }), .B_DOUT({nc1245, nc1246, nc1247, 
        nc1248, nc1249, nc1250, nc1251, nc1252, nc1253, nc1254, nc1255, 
        nc1256, nc1257, nc1258, nc1259, \B_DOUT_TEMPR68[34] , 
        \B_DOUT_TEMPR68[33] , \B_DOUT_TEMPR68[32] , 
        \B_DOUT_TEMPR68[31] , \B_DOUT_TEMPR68[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[68][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%113%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R113C2 (
        .A_DOUT({nc1260, nc1261, nc1262, nc1263, nc1264, nc1265, 
        nc1266, nc1267, nc1268, nc1269, nc1270, nc1271, nc1272, nc1273, 
        nc1274, \A_DOUT_TEMPR113[14] , \A_DOUT_TEMPR113[13] , 
        \A_DOUT_TEMPR113[12] , \A_DOUT_TEMPR113[11] , 
        \A_DOUT_TEMPR113[10] }), .B_DOUT({nc1275, nc1276, nc1277, 
        nc1278, nc1279, nc1280, nc1281, nc1282, nc1283, nc1284, nc1285, 
        nc1286, nc1287, nc1288, nc1289, \B_DOUT_TEMPR113[14] , 
        \B_DOUT_TEMPR113[13] , \B_DOUT_TEMPR113[12] , 
        \B_DOUT_TEMPR113[11] , \B_DOUT_TEMPR113[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[113][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_3036 (.A(\A_DOUT_TEMPR99[24] ), .B(\A_DOUT_TEMPR100[24] ), 
        .C(\A_DOUT_TEMPR101[24] ), .D(\A_DOUT_TEMPR102[24] ), .Y(
        OR4_3036_Y));
    OR4 OR4_1967 (.A(\A_DOUT_TEMPR28[36] ), .B(\A_DOUT_TEMPR29[36] ), 
        .C(\A_DOUT_TEMPR30[36] ), .D(\A_DOUT_TEMPR31[36] ), .Y(
        OR4_1967_Y));
    OR4 OR4_360 (.A(OR4_1533_Y), .B(OR4_1925_Y), .C(OR4_2678_Y), .D(
        OR4_434_Y), .Y(OR4_360_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%52%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R52C6 (
        .A_DOUT({nc1290, nc1291, nc1292, nc1293, nc1294, nc1295, 
        nc1296, nc1297, nc1298, nc1299, nc1300, nc1301, nc1302, nc1303, 
        nc1304, \A_DOUT_TEMPR52[34] , \A_DOUT_TEMPR52[33] , 
        \A_DOUT_TEMPR52[32] , \A_DOUT_TEMPR52[31] , 
        \A_DOUT_TEMPR52[30] }), .B_DOUT({nc1305, nc1306, nc1307, 
        nc1308, nc1309, nc1310, nc1311, nc1312, nc1313, nc1314, nc1315, 
        nc1316, nc1317, nc1318, nc1319, \B_DOUT_TEMPR52[34] , 
        \B_DOUT_TEMPR52[33] , \B_DOUT_TEMPR52[32] , 
        \B_DOUT_TEMPR52[31] , \B_DOUT_TEMPR52[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[52][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1208 (.A(\A_DOUT_TEMPR0[6] ), .B(\A_DOUT_TEMPR1[6] ), .C(
        \A_DOUT_TEMPR2[6] ), .D(\A_DOUT_TEMPR3[6] ), .Y(OR4_1208_Y));
    OR4 OR4_1318 (.A(\B_DOUT_TEMPR60[4] ), .B(\B_DOUT_TEMPR61[4] ), .C(
        \B_DOUT_TEMPR62[4] ), .D(\B_DOUT_TEMPR63[4] ), .Y(OR4_1318_Y));
    OR4 OR4_347 (.A(OR4_1185_Y), .B(OR4_338_Y), .C(OR4_2353_Y), .D(
        OR4_2679_Y), .Y(OR4_347_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%59%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R59C0 (
        .A_DOUT({nc1320, nc1321, nc1322, nc1323, nc1324, nc1325, 
        nc1326, nc1327, nc1328, nc1329, nc1330, nc1331, nc1332, nc1333, 
        nc1334, \A_DOUT_TEMPR59[4] , \A_DOUT_TEMPR59[3] , 
        \A_DOUT_TEMPR59[2] , \A_DOUT_TEMPR59[1] , \A_DOUT_TEMPR59[0] })
        , .B_DOUT({nc1335, nc1336, nc1337, nc1338, nc1339, nc1340, 
        nc1341, nc1342, nc1343, nc1344, nc1345, nc1346, nc1347, nc1348, 
        nc1349, \B_DOUT_TEMPR59[4] , \B_DOUT_TEMPR59[3] , 
        \B_DOUT_TEMPR59[2] , \B_DOUT_TEMPR59[1] , \B_DOUT_TEMPR59[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[59][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2275 (.A(\B_DOUT_TEMPR91[23] ), .B(\B_DOUT_TEMPR92[23] ), 
        .C(\B_DOUT_TEMPR93[23] ), .D(\B_DOUT_TEMPR94[23] ), .Y(
        OR4_2275_Y));
    OR4 OR4_1450 (.A(\B_DOUT_TEMPR12[27] ), .B(\B_DOUT_TEMPR13[27] ), 
        .C(\B_DOUT_TEMPR14[27] ), .D(\B_DOUT_TEMPR15[27] ), .Y(
        OR4_1450_Y));
    OR4 OR4_848 (.A(\B_DOUT_TEMPR83[35] ), .B(\B_DOUT_TEMPR84[35] ), 
        .C(\B_DOUT_TEMPR85[35] ), .D(\B_DOUT_TEMPR86[35] ), .Y(
        OR4_848_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%95%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R95C2 (
        .A_DOUT({nc1350, nc1351, nc1352, nc1353, nc1354, nc1355, 
        nc1356, nc1357, nc1358, nc1359, nc1360, nc1361, nc1362, nc1363, 
        nc1364, \A_DOUT_TEMPR95[14] , \A_DOUT_TEMPR95[13] , 
        \A_DOUT_TEMPR95[12] , \A_DOUT_TEMPR95[11] , 
        \A_DOUT_TEMPR95[10] }), .B_DOUT({nc1365, nc1366, nc1367, 
        nc1368, nc1369, nc1370, nc1371, nc1372, nc1373, nc1374, nc1375, 
        nc1376, nc1377, nc1378, nc1379, \B_DOUT_TEMPR95[14] , 
        \B_DOUT_TEMPR95[13] , \B_DOUT_TEMPR95[12] , 
        \B_DOUT_TEMPR95[11] , \B_DOUT_TEMPR95[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[95][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1283 (.A(\A_DOUT_TEMPR111[36] ), .B(\A_DOUT_TEMPR112[36] ), 
        .C(\A_DOUT_TEMPR113[36] ), .D(\A_DOUT_TEMPR114[36] ), .Y(
        OR4_1283_Y));
    OR4 OR4_1974 (.A(OR4_226_Y), .B(OR4_1299_Y), .C(OR4_2999_Y), .D(
        OR4_1383_Y), .Y(OR4_1974_Y));
    OR4 OR4_641 (.A(OR4_1053_Y), .B(OR4_2743_Y), .C(OR4_1068_Y), .D(
        OR4_1347_Y), .Y(OR4_641_Y));
    OR4 OR4_2663 (.A(\A_DOUT_TEMPR99[2] ), .B(\A_DOUT_TEMPR100[2] ), 
        .C(\A_DOUT_TEMPR101[2] ), .D(\A_DOUT_TEMPR102[2] ), .Y(
        OR4_2663_Y));
    OR4 OR4_2921 (.A(OR4_1063_Y), .B(OR4_2456_Y), .C(OR2_48_Y), .D(
        \A_DOUT_TEMPR74[5] ), .Y(OR4_2921_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%55%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R55C6 (
        .A_DOUT({nc1380, nc1381, nc1382, nc1383, nc1384, nc1385, 
        nc1386, nc1387, nc1388, nc1389, nc1390, nc1391, nc1392, nc1393, 
        nc1394, \A_DOUT_TEMPR55[34] , \A_DOUT_TEMPR55[33] , 
        \A_DOUT_TEMPR55[32] , \A_DOUT_TEMPR55[31] , 
        \A_DOUT_TEMPR55[30] }), .B_DOUT({nc1395, nc1396, nc1397, 
        nc1398, nc1399, nc1400, nc1401, nc1402, nc1403, nc1404, nc1405, 
        nc1406, nc1407, nc1408, nc1409, \B_DOUT_TEMPR55[34] , 
        \B_DOUT_TEMPR55[33] , \B_DOUT_TEMPR55[32] , 
        \B_DOUT_TEMPR55[31] , \B_DOUT_TEMPR55[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[55][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2969 (.A(\A_DOUT_TEMPR95[18] ), .B(\A_DOUT_TEMPR96[18] ), 
        .C(\A_DOUT_TEMPR97[18] ), .D(\A_DOUT_TEMPR98[18] ), .Y(
        OR4_2969_Y));
    OR4 OR4_1860 (.A(\B_DOUT_TEMPR60[29] ), .B(\B_DOUT_TEMPR61[29] ), 
        .C(\B_DOUT_TEMPR62[29] ), .D(\B_DOUT_TEMPR63[29] ), .Y(
        OR4_1860_Y));
    OR4 OR4_1976 (.A(\B_DOUT_TEMPR20[24] ), .B(\B_DOUT_TEMPR21[24] ), 
        .C(\B_DOUT_TEMPR22[24] ), .D(\B_DOUT_TEMPR23[24] ), .Y(
        OR4_1976_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%10%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R10C0 (
        .A_DOUT({nc1410, nc1411, nc1412, nc1413, nc1414, nc1415, 
        nc1416, nc1417, nc1418, nc1419, nc1420, nc1421, nc1422, nc1423, 
        nc1424, \A_DOUT_TEMPR10[4] , \A_DOUT_TEMPR10[3] , 
        \A_DOUT_TEMPR10[2] , \A_DOUT_TEMPR10[1] , \A_DOUT_TEMPR10[0] })
        , .B_DOUT({nc1425, nc1426, nc1427, nc1428, nc1429, nc1430, 
        nc1431, nc1432, nc1433, nc1434, nc1435, nc1436, nc1437, nc1438, 
        nc1439, \B_DOUT_TEMPR10[4] , \B_DOUT_TEMPR10[3] , 
        \B_DOUT_TEMPR10[2] , \B_DOUT_TEMPR10[1] , \B_DOUT_TEMPR10[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[10][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_44 (.A(\A_DOUT_TEMPR28[33] ), .B(\A_DOUT_TEMPR29[33] ), .C(
        \A_DOUT_TEMPR30[33] ), .D(\A_DOUT_TEMPR31[33] ), .Y(OR4_44_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%15%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R15C4 (
        .A_DOUT({nc1440, nc1441, nc1442, nc1443, nc1444, nc1445, 
        nc1446, nc1447, nc1448, nc1449, nc1450, nc1451, nc1452, nc1453, 
        nc1454, \A_DOUT_TEMPR15[24] , \A_DOUT_TEMPR15[23] , 
        \A_DOUT_TEMPR15[22] , \A_DOUT_TEMPR15[21] , 
        \A_DOUT_TEMPR15[20] }), .B_DOUT({nc1455, nc1456, nc1457, 
        nc1458, nc1459, nc1460, nc1461, nc1462, nc1463, nc1464, nc1465, 
        nc1466, nc1467, nc1468, nc1469, \B_DOUT_TEMPR15[24] , 
        \B_DOUT_TEMPR15[23] , \B_DOUT_TEMPR15[22] , 
        \B_DOUT_TEMPR15[21] , \B_DOUT_TEMPR15[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[15][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1255 (.A(\A_DOUT_TEMPR4[28] ), .B(\A_DOUT_TEMPR5[28] ), .C(
        \A_DOUT_TEMPR6[28] ), .D(\A_DOUT_TEMPR7[28] ), .Y(OR4_1255_Y));
    OR4 OR4_444 (.A(OR4_1897_Y), .B(OR4_1102_Y), .C(OR4_662_Y), .D(
        OR4_2315_Y), .Y(OR4_444_Y));
    OR4 OR4_2358 (.A(\B_DOUT_TEMPR68[14] ), .B(\B_DOUT_TEMPR69[14] ), 
        .C(\B_DOUT_TEMPR70[14] ), .D(\B_DOUT_TEMPR71[14] ), .Y(
        OR4_2358_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%64%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R64C3 (
        .A_DOUT({nc1470, nc1471, nc1472, nc1473, nc1474, nc1475, 
        nc1476, nc1477, nc1478, nc1479, nc1480, nc1481, nc1482, nc1483, 
        nc1484, \A_DOUT_TEMPR64[19] , \A_DOUT_TEMPR64[18] , 
        \A_DOUT_TEMPR64[17] , \A_DOUT_TEMPR64[16] , 
        \A_DOUT_TEMPR64[15] }), .B_DOUT({nc1485, nc1486, nc1487, 
        nc1488, nc1489, nc1490, nc1491, nc1492, nc1493, nc1494, nc1495, 
        nc1496, nc1497, nc1498, nc1499, \B_DOUT_TEMPR64[19] , 
        \B_DOUT_TEMPR64[18] , \B_DOUT_TEMPR64[17] , 
        \B_DOUT_TEMPR64[16] , \B_DOUT_TEMPR64[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[64][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1864 (.A(\B_DOUT_TEMPR44[35] ), .B(\B_DOUT_TEMPR45[35] ), 
        .C(\B_DOUT_TEMPR46[35] ), .D(\B_DOUT_TEMPR47[35] ), .Y(
        OR4_1864_Y));
    OR4 OR4_1198 (.A(\A_DOUT_TEMPR83[1] ), .B(\A_DOUT_TEMPR84[1] ), .C(
        \A_DOUT_TEMPR85[1] ), .D(\A_DOUT_TEMPR86[1] ), .Y(OR4_1198_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%5%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R5C7 (
        .A_DOUT({nc1500, nc1501, nc1502, nc1503, nc1504, nc1505, 
        nc1506, nc1507, nc1508, nc1509, nc1510, nc1511, nc1512, nc1513, 
        nc1514, \A_DOUT_TEMPR5[39] , \A_DOUT_TEMPR5[38] , 
        \A_DOUT_TEMPR5[37] , \A_DOUT_TEMPR5[36] , \A_DOUT_TEMPR5[35] })
        , .B_DOUT({nc1515, nc1516, nc1517, nc1518, nc1519, nc1520, 
        nc1521, nc1522, nc1523, nc1524, nc1525, nc1526, nc1527, nc1528, 
        nc1529, \B_DOUT_TEMPR5[39] , \B_DOUT_TEMPR5[38] , 
        \B_DOUT_TEMPR5[37] , \B_DOUT_TEMPR5[36] , \B_DOUT_TEMPR5[35] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[5][7] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[39], A_DIN[38], A_DIN[37], 
        A_DIN[36], A_DIN[35]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_430 (.A(\B_DOUT_TEMPR75[4] ), .B(\B_DOUT_TEMPR76[4] ), .C(
        \B_DOUT_TEMPR77[4] ), .D(\B_DOUT_TEMPR78[4] ), .Y(OR4_430_Y));
    OR4 OR4_290 (.A(\B_DOUT_TEMPR52[14] ), .B(\B_DOUT_TEMPR53[14] ), 
        .C(\B_DOUT_TEMPR54[14] ), .D(\B_DOUT_TEMPR55[14] ), .Y(
        OR4_290_Y));
    OR4 OR4_2200 (.A(OR4_650_Y), .B(OR4_1099_Y), .C(OR4_261_Y), .D(
        OR4_2213_Y), .Y(OR4_2200_Y));
    OR4 OR4_2838 (.A(\B_DOUT_TEMPR56[13] ), .B(\B_DOUT_TEMPR57[13] ), 
        .C(\B_DOUT_TEMPR58[13] ), .D(\B_DOUT_TEMPR59[13] ), .Y(
        OR4_2838_Y));
    OR4 OR4_2764 (.A(\A_DOUT_TEMPR107[2] ), .B(\A_DOUT_TEMPR108[2] ), 
        .C(\A_DOUT_TEMPR109[2] ), .D(\A_DOUT_TEMPR110[2] ), .Y(
        OR4_2764_Y));
    OR4 OR4_690 (.A(OR4_2295_Y), .B(OR4_2619_Y), .C(OR4_2218_Y), .D(
        OR4_2638_Y), .Y(OR4_690_Y));
    OR4 OR4_3002 (.A(\A_DOUT_TEMPR32[22] ), .B(\A_DOUT_TEMPR33[22] ), 
        .C(\A_DOUT_TEMPR34[22] ), .D(\A_DOUT_TEMPR35[22] ), .Y(
        OR4_3002_Y));
    OR4 OR4_824 (.A(OR4_1330_Y), .B(OR4_1260_Y), .C(OR4_1942_Y), .D(
        OR4_2209_Y), .Y(OR4_824_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[0]  (.A(CFG3_11_Y), .B(
        CFG3_16_Y), .Y(\BLKY2[0] ));
    OR4 OR4_2461 (.A(\B_DOUT_TEMPR56[16] ), .B(\B_DOUT_TEMPR57[16] ), 
        .C(\B_DOUT_TEMPR58[16] ), .D(\B_DOUT_TEMPR59[16] ), .Y(
        OR4_2461_Y));
    OR4 OR4_1838 (.A(\A_DOUT_TEMPR64[20] ), .B(\A_DOUT_TEMPR65[20] ), 
        .C(\A_DOUT_TEMPR66[20] ), .D(\A_DOUT_TEMPR67[20] ), .Y(
        OR4_1838_Y));
    OR4 OR4_1415 (.A(\B_DOUT_TEMPR24[30] ), .B(\B_DOUT_TEMPR25[30] ), 
        .C(\B_DOUT_TEMPR26[30] ), .D(\B_DOUT_TEMPR27[30] ), .Y(
        OR4_1415_Y));
    OR4 OR4_522 (.A(OR4_472_Y), .B(OR4_766_Y), .C(OR4_401_Y), .D(
        OR4_782_Y), .Y(OR4_522_Y));
    OR4 OR4_2223 (.A(\B_DOUT_TEMPR56[5] ), .B(\B_DOUT_TEMPR57[5] ), .C(
        \B_DOUT_TEMPR58[5] ), .D(\B_DOUT_TEMPR59[5] ), .Y(OR4_2223_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%32%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R32C6 (
        .A_DOUT({nc1530, nc1531, nc1532, nc1533, nc1534, nc1535, 
        nc1536, nc1537, nc1538, nc1539, nc1540, nc1541, nc1542, nc1543, 
        nc1544, \A_DOUT_TEMPR32[34] , \A_DOUT_TEMPR32[33] , 
        \A_DOUT_TEMPR32[32] , \A_DOUT_TEMPR32[31] , 
        \A_DOUT_TEMPR32[30] }), .B_DOUT({nc1545, nc1546, nc1547, 
        nc1548, nc1549, nc1550, nc1551, nc1552, nc1553, nc1554, nc1555, 
        nc1556, nc1557, nc1558, nc1559, \B_DOUT_TEMPR32[34] , 
        \B_DOUT_TEMPR32[33] , \B_DOUT_TEMPR32[32] , 
        \B_DOUT_TEMPR32[31] , \B_DOUT_TEMPR32[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[32][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_17 (.A(\B_DOUT_TEMPR111[7] ), .B(\B_DOUT_TEMPR112[7] ), .C(
        \B_DOUT_TEMPR113[7] ), .D(\B_DOUT_TEMPR114[7] ), .Y(OR4_17_Y));
    OR4 OR4_779 (.A(\A_DOUT_TEMPR44[16] ), .B(\A_DOUT_TEMPR45[16] ), 
        .C(\A_DOUT_TEMPR46[16] ), .D(\A_DOUT_TEMPR47[16] ), .Y(
        OR4_779_Y));
    OR4 OR4_1893 (.A(\A_DOUT_TEMPR0[34] ), .B(\A_DOUT_TEMPR1[34] ), .C(
        \A_DOUT_TEMPR2[34] ), .D(\A_DOUT_TEMPR3[34] ), .Y(OR4_1893_Y));
    OR2 OR2_2 (.A(\B_DOUT_TEMPR72[9] ), .B(\B_DOUT_TEMPR73[9] ), .Y(
        OR2_2_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%78%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R78C1 (
        .A_DOUT({nc1560, nc1561, nc1562, nc1563, nc1564, nc1565, 
        nc1566, nc1567, nc1568, nc1569, nc1570, nc1571, nc1572, nc1573, 
        nc1574, \A_DOUT_TEMPR78[9] , \A_DOUT_TEMPR78[8] , 
        \A_DOUT_TEMPR78[7] , \A_DOUT_TEMPR78[6] , \A_DOUT_TEMPR78[5] })
        , .B_DOUT({nc1575, nc1576, nc1577, nc1578, nc1579, nc1580, 
        nc1581, nc1582, nc1583, nc1584, nc1585, nc1586, nc1587, nc1588, 
        nc1589, \B_DOUT_TEMPR78[9] , \B_DOUT_TEMPR78[8] , 
        \B_DOUT_TEMPR78[7] , \B_DOUT_TEMPR78[6] , \B_DOUT_TEMPR78[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[78][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[18]  (.A(OR4_30_Y), .B(OR4_2326_Y), .C(OR4_1755_Y), 
        .D(OR4_2164_Y), .Y(A_DOUT[18]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%39%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R39C0 (
        .A_DOUT({nc1590, nc1591, nc1592, nc1593, nc1594, nc1595, 
        nc1596, nc1597, nc1598, nc1599, nc1600, nc1601, nc1602, nc1603, 
        nc1604, \A_DOUT_TEMPR39[4] , \A_DOUT_TEMPR39[3] , 
        \A_DOUT_TEMPR39[2] , \A_DOUT_TEMPR39[1] , \A_DOUT_TEMPR39[0] })
        , .B_DOUT({nc1605, nc1606, nc1607, nc1608, nc1609, nc1610, 
        nc1611, nc1612, nc1613, nc1614, nc1615, nc1616, nc1617, nc1618, 
        nc1619, \B_DOUT_TEMPR39[4] , \B_DOUT_TEMPR39[3] , 
        \B_DOUT_TEMPR39[2] , \B_DOUT_TEMPR39[1] , \B_DOUT_TEMPR39[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[39][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%78%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R78C7 (
        .A_DOUT({nc1620, nc1621, nc1622, nc1623, nc1624, nc1625, 
        nc1626, nc1627, nc1628, nc1629, nc1630, nc1631, nc1632, nc1633, 
        nc1634, \A_DOUT_TEMPR78[39] , \A_DOUT_TEMPR78[38] , 
        \A_DOUT_TEMPR78[37] , \A_DOUT_TEMPR78[36] , 
        \A_DOUT_TEMPR78[35] }), .B_DOUT({nc1635, nc1636, nc1637, 
        nc1638, nc1639, nc1640, nc1641, nc1642, nc1643, nc1644, nc1645, 
        nc1646, nc1647, nc1648, nc1649, \B_DOUT_TEMPR78[39] , 
        \B_DOUT_TEMPR78[38] , \B_DOUT_TEMPR78[37] , 
        \B_DOUT_TEMPR78[36] , \B_DOUT_TEMPR78[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[78][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_675 (.A(OR4_1470_Y), .B(OR4_791_Y), .C(OR4_1480_Y), .D(
        OR4_1775_Y), .Y(OR4_675_Y));
    OR4 OR4_1799 (.A(\B_DOUT_TEMPR12[5] ), .B(\B_DOUT_TEMPR13[5] ), .C(
        \B_DOUT_TEMPR14[5] ), .D(\B_DOUT_TEMPR15[5] ), .Y(OR4_1799_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%102%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R102C2 (
        .A_DOUT({nc1650, nc1651, nc1652, nc1653, nc1654, nc1655, 
        nc1656, nc1657, nc1658, nc1659, nc1660, nc1661, nc1662, nc1663, 
        nc1664, \A_DOUT_TEMPR102[14] , \A_DOUT_TEMPR102[13] , 
        \A_DOUT_TEMPR102[12] , \A_DOUT_TEMPR102[11] , 
        \A_DOUT_TEMPR102[10] }), .B_DOUT({nc1665, nc1666, nc1667, 
        nc1668, nc1669, nc1670, nc1671, nc1672, nc1673, nc1674, nc1675, 
        nc1676, nc1677, nc1678, nc1679, \B_DOUT_TEMPR102[14] , 
        \B_DOUT_TEMPR102[13] , \B_DOUT_TEMPR102[12] , 
        \B_DOUT_TEMPR102[11] , \B_DOUT_TEMPR102[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[102][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_264 (.A(OR4_1703_Y), .B(OR4_1528_Y), .C(OR2_34_Y), .D(
        \A_DOUT_TEMPR74[38] ), .Y(OR4_264_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[14]  (.A(CFG3_0_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[14] ));
    OR4 OR4_2306 (.A(OR4_1192_Y), .B(OR4_1966_Y), .C(OR4_2675_Y), .D(
        OR4_2973_Y), .Y(OR4_2306_Y));
    OR4 OR4_279 (.A(\A_DOUT_TEMPR36[27] ), .B(\A_DOUT_TEMPR37[27] ), 
        .C(\A_DOUT_TEMPR38[27] ), .D(\A_DOUT_TEMPR39[27] ), .Y(
        OR4_279_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%111%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R111C5 (
        .A_DOUT({nc1680, nc1681, nc1682, nc1683, nc1684, nc1685, 
        nc1686, nc1687, nc1688, nc1689, nc1690, nc1691, nc1692, nc1693, 
        nc1694, \A_DOUT_TEMPR111[29] , \A_DOUT_TEMPR111[28] , 
        \A_DOUT_TEMPR111[27] , \A_DOUT_TEMPR111[26] , 
        \A_DOUT_TEMPR111[25] }), .B_DOUT({nc1695, nc1696, nc1697, 
        nc1698, nc1699, nc1700, nc1701, nc1702, nc1703, nc1704, nc1705, 
        nc1706, nc1707, nc1708, nc1709, \B_DOUT_TEMPR111[29] , 
        \B_DOUT_TEMPR111[28] , \B_DOUT_TEMPR111[27] , 
        \B_DOUT_TEMPR111[26] , \B_DOUT_TEMPR111[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[111][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2618 (.A(\A_DOUT_TEMPR60[10] ), .B(\A_DOUT_TEMPR61[10] ), 
        .C(\A_DOUT_TEMPR62[10] ), .D(\A_DOUT_TEMPR63[10] ), .Y(
        OR4_2618_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%35%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R35C6 (
        .A_DOUT({nc1710, nc1711, nc1712, nc1713, nc1714, nc1715, 
        nc1716, nc1717, nc1718, nc1719, nc1720, nc1721, nc1722, nc1723, 
        nc1724, \A_DOUT_TEMPR35[34] , \A_DOUT_TEMPR35[33] , 
        \A_DOUT_TEMPR35[32] , \A_DOUT_TEMPR35[31] , 
        \A_DOUT_TEMPR35[30] }), .B_DOUT({nc1725, nc1726, nc1727, 
        nc1728, nc1729, nc1730, nc1731, nc1732, nc1733, nc1734, nc1735, 
        nc1736, nc1737, nc1738, nc1739, \B_DOUT_TEMPR35[34] , 
        \B_DOUT_TEMPR35[33] , \B_DOUT_TEMPR35[32] , 
        \B_DOUT_TEMPR35[31] , \B_DOUT_TEMPR35[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[35][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%86%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R86C0 (
        .A_DOUT({nc1740, nc1741, nc1742, nc1743, nc1744, nc1745, 
        nc1746, nc1747, nc1748, nc1749, nc1750, nc1751, nc1752, nc1753, 
        nc1754, \A_DOUT_TEMPR86[4] , \A_DOUT_TEMPR86[3] , 
        \A_DOUT_TEMPR86[2] , \A_DOUT_TEMPR86[1] , \A_DOUT_TEMPR86[0] })
        , .B_DOUT({nc1755, nc1756, nc1757, nc1758, nc1759, nc1760, 
        nc1761, nc1762, nc1763, nc1764, nc1765, nc1766, nc1767, nc1768, 
        nc1769, \B_DOUT_TEMPR86[4] , \B_DOUT_TEMPR86[3] , 
        \B_DOUT_TEMPR86[2] , \B_DOUT_TEMPR86[1] , \B_DOUT_TEMPR86[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[86][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_760 (.A(\B_DOUT_TEMPR0[35] ), .B(\B_DOUT_TEMPR1[35] ), .C(
        \B_DOUT_TEMPR2[35] ), .D(\B_DOUT_TEMPR3[35] ), .Y(OR4_760_Y));
    OR4 OR4_2676 (.A(\B_DOUT_TEMPR20[37] ), .B(\B_DOUT_TEMPR21[37] ), 
        .C(\B_DOUT_TEMPR22[37] ), .D(\B_DOUT_TEMPR23[37] ), .Y(
        OR4_2676_Y));
    OR4 OR4_773 (.A(\A_DOUT_TEMPR99[39] ), .B(\A_DOUT_TEMPR100[39] ), 
        .C(\A_DOUT_TEMPR101[39] ), .D(\A_DOUT_TEMPR102[39] ), .Y(
        OR4_773_Y));
    OR4 OR4_1716 (.A(OR4_1079_Y), .B(OR4_2785_Y), .C(OR4_344_Y), .D(
        OR4_2592_Y), .Y(OR4_1716_Y));
    OR4 OR4_1196 (.A(\B_DOUT_TEMPR91[32] ), .B(\B_DOUT_TEMPR92[32] ), 
        .C(\B_DOUT_TEMPR93[32] ), .D(\B_DOUT_TEMPR94[32] ), .Y(
        OR4_1196_Y));
    OR4 OR4_2170 (.A(\B_DOUT_TEMPR36[25] ), .B(\B_DOUT_TEMPR37[25] ), 
        .C(\B_DOUT_TEMPR38[25] ), .D(\B_DOUT_TEMPR39[25] ), .Y(
        OR4_2170_Y));
    OR4 OR4_2455 (.A(\A_DOUT_TEMPR95[12] ), .B(\A_DOUT_TEMPR96[12] ), 
        .C(\A_DOUT_TEMPR97[12] ), .D(\A_DOUT_TEMPR98[12] ), .Y(
        OR4_2455_Y));
    OR4 OR4_1598 (.A(\A_DOUT_TEMPR52[15] ), .B(\A_DOUT_TEMPR53[15] ), 
        .C(\A_DOUT_TEMPR54[15] ), .D(\A_DOUT_TEMPR55[15] ), .Y(
        OR4_1598_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%112%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R112C0 (
        .A_DOUT({nc1770, nc1771, nc1772, nc1773, nc1774, nc1775, 
        nc1776, nc1777, nc1778, nc1779, nc1780, nc1781, nc1782, nc1783, 
        nc1784, \A_DOUT_TEMPR112[4] , \A_DOUT_TEMPR112[3] , 
        \A_DOUT_TEMPR112[2] , \A_DOUT_TEMPR112[1] , 
        \A_DOUT_TEMPR112[0] }), .B_DOUT({nc1785, nc1786, nc1787, 
        nc1788, nc1789, nc1790, nc1791, nc1792, nc1793, nc1794, nc1795, 
        nc1796, nc1797, nc1798, nc1799, \B_DOUT_TEMPR112[4] , 
        \B_DOUT_TEMPR112[3] , \B_DOUT_TEMPR112[2] , 
        \B_DOUT_TEMPR112[1] , \B_DOUT_TEMPR112[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[112][0] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[4], 
        B_DIN[3], B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_139 (.A(\A_DOUT_TEMPR83[39] ), .B(\A_DOUT_TEMPR84[39] ), 
        .C(\A_DOUT_TEMPR85[39] ), .D(\A_DOUT_TEMPR86[39] ), .Y(
        OR4_139_Y));
    OR4 OR4_2964 (.A(\B_DOUT_TEMPR91[24] ), .B(\B_DOUT_TEMPR92[24] ), 
        .C(\B_DOUT_TEMPR93[24] ), .D(\B_DOUT_TEMPR94[24] ), .Y(
        OR4_2964_Y));
    OR4 OR4_1348 (.A(\A_DOUT_TEMPR95[21] ), .B(\A_DOUT_TEMPR96[21] ), 
        .C(\A_DOUT_TEMPR97[21] ), .D(\A_DOUT_TEMPR98[21] ), .Y(
        OR4_1348_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[27]  (.A(CFG3_23_Y), .B(
        CFG3_18_Y), .Y(\BLKX2[27] ));
    OR4 OR4_2738 (.A(\A_DOUT_TEMPR95[34] ), .B(\A_DOUT_TEMPR96[34] ), 
        .C(\A_DOUT_TEMPR97[34] ), .D(\A_DOUT_TEMPR98[34] ), .Y(
        OR4_2738_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%18%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R18C6 (
        .A_DOUT({nc1800, nc1801, nc1802, nc1803, nc1804, nc1805, 
        nc1806, nc1807, nc1808, nc1809, nc1810, nc1811, nc1812, nc1813, 
        nc1814, \A_DOUT_TEMPR18[34] , \A_DOUT_TEMPR18[33] , 
        \A_DOUT_TEMPR18[32] , \A_DOUT_TEMPR18[31] , 
        \A_DOUT_TEMPR18[30] }), .B_DOUT({nc1815, nc1816, nc1817, 
        nc1818, nc1819, nc1820, nc1821, nc1822, nc1823, nc1824, nc1825, 
        nc1826, nc1827, nc1828, nc1829, \B_DOUT_TEMPR18[34] , 
        \B_DOUT_TEMPR18[33] , \B_DOUT_TEMPR18[32] , 
        \B_DOUT_TEMPR18[31] , \B_DOUT_TEMPR18[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[18][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2966 (.A(\A_DOUT_TEMPR115[11] ), .B(\A_DOUT_TEMPR116[11] ), 
        .C(\A_DOUT_TEMPR117[11] ), .D(\A_DOUT_TEMPR118[11] ), .Y(
        OR4_2966_Y));
    OR4 OR4_278 (.A(\B_DOUT_TEMPR95[3] ), .B(\B_DOUT_TEMPR96[3] ), .C(
        \B_DOUT_TEMPR97[3] ), .D(\B_DOUT_TEMPR98[3] ), .Y(OR4_278_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%115%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R115C1 (
        .A_DOUT({nc1830, nc1831, nc1832, nc1833, nc1834, nc1835, 
        nc1836, nc1837, nc1838, nc1839, nc1840, nc1841, nc1842, nc1843, 
        nc1844, \A_DOUT_TEMPR115[9] , \A_DOUT_TEMPR115[8] , 
        \A_DOUT_TEMPR115[7] , \A_DOUT_TEMPR115[6] , 
        \A_DOUT_TEMPR115[5] }), .B_DOUT({nc1845, nc1846, nc1847, 
        nc1848, nc1849, nc1850, nc1851, nc1852, nc1853, nc1854, nc1855, 
        nc1856, nc1857, nc1858, nc1859, \B_DOUT_TEMPR115[9] , 
        \B_DOUT_TEMPR115[8] , \B_DOUT_TEMPR115[7] , 
        \B_DOUT_TEMPR115[6] , \B_DOUT_TEMPR115[5] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[115][1] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[9], 
        B_DIN[8], B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1024 (.A(OR4_801_Y), .B(OR4_1704_Y), .C(OR4_1376_Y), .D(
        OR4_2884_Y), .Y(OR4_1024_Y));
    OR4 OR4_1026 (.A(\B_DOUT_TEMPR87[39] ), .B(\B_DOUT_TEMPR88[39] ), 
        .C(\B_DOUT_TEMPR89[39] ), .D(\B_DOUT_TEMPR90[39] ), .Y(
        OR4_1026_Y));
    OR4 OR4_1656 (.A(\B_DOUT_TEMPR64[8] ), .B(\B_DOUT_TEMPR65[8] ), .C(
        \B_DOUT_TEMPR66[8] ), .D(\B_DOUT_TEMPR67[8] ), .Y(OR4_1656_Y));
    OR4 OR4_10 (.A(\B_DOUT_TEMPR28[27] ), .B(\B_DOUT_TEMPR29[27] ), .C(
        \B_DOUT_TEMPR30[27] ), .D(\B_DOUT_TEMPR31[27] ), .Y(OR4_10_Y));
    OR4 OR4_709 (.A(\B_DOUT_TEMPR24[34] ), .B(\B_DOUT_TEMPR25[34] ), 
        .C(\B_DOUT_TEMPR26[34] ), .D(\B_DOUT_TEMPR27[34] ), .Y(
        OR4_709_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKY0[0]  (.A(B_ADDR[12]), .Y(
        \BLKY0[0] ));
    OR4 OR4_1738 (.A(\A_DOUT_TEMPR56[4] ), .B(\A_DOUT_TEMPR57[4] ), .C(
        \A_DOUT_TEMPR58[4] ), .D(\A_DOUT_TEMPR59[4] ), .Y(OR4_1738_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%92%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R92C5 (
        .A_DOUT({nc1860, nc1861, nc1862, nc1863, nc1864, nc1865, 
        nc1866, nc1867, nc1868, nc1869, nc1870, nc1871, nc1872, nc1873, 
        nc1874, \A_DOUT_TEMPR92[29] , \A_DOUT_TEMPR92[28] , 
        \A_DOUT_TEMPR92[27] , \A_DOUT_TEMPR92[26] , 
        \A_DOUT_TEMPR92[25] }), .B_DOUT({nc1875, nc1876, nc1877, 
        nc1878, nc1879, nc1880, nc1881, nc1882, nc1883, nc1884, nc1885, 
        nc1886, nc1887, nc1888, nc1889, \B_DOUT_TEMPR92[29] , 
        \B_DOUT_TEMPR92[28] , \B_DOUT_TEMPR92[27] , 
        \B_DOUT_TEMPR92[26] , \B_DOUT_TEMPR92[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[92][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2543 (.A(\A_DOUT_TEMPR79[1] ), .B(\A_DOUT_TEMPR80[1] ), .C(
        \A_DOUT_TEMPR81[1] ), .D(\A_DOUT_TEMPR82[1] ), .Y(OR4_2543_Y));
    OR4 OR4_1150 (.A(OR4_1602_Y), .B(OR4_787_Y), .C(OR4_2826_Y), .D(
        OR4_67_Y), .Y(OR4_1150_Y));
    OR4 OR4_844 (.A(OR4_2978_Y), .B(OR4_1899_Y), .C(OR4_520_Y), .D(
        OR4_1499_Y), .Y(OR4_844_Y));
    OR4 OR4_605 (.A(OR4_497_Y), .B(OR4_1798_Y), .C(OR4_2430_Y), .D(
        OR4_1617_Y), .Y(OR4_605_Y));
    OR4 OR4_2143 (.A(\A_DOUT_TEMPR24[36] ), .B(\A_DOUT_TEMPR25[36] ), 
        .C(\A_DOUT_TEMPR26[36] ), .D(\A_DOUT_TEMPR27[36] ), .Y(
        OR4_2143_Y));
    OR4 OR4_2756 (.A(\A_DOUT_TEMPR44[39] ), .B(\A_DOUT_TEMPR45[39] ), 
        .C(\A_DOUT_TEMPR46[39] ), .D(\A_DOUT_TEMPR47[39] ), .Y(
        OR4_2756_Y));
    OR4 OR4_542 (.A(\B_DOUT_TEMPR79[35] ), .B(\B_DOUT_TEMPR80[35] ), 
        .C(\B_DOUT_TEMPR81[35] ), .D(\B_DOUT_TEMPR82[35] ), .Y(
        OR4_542_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%71%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R71C1 (
        .A_DOUT({nc1890, nc1891, nc1892, nc1893, nc1894, nc1895, 
        nc1896, nc1897, nc1898, nc1899, nc1900, nc1901, nc1902, nc1903, 
        nc1904, \A_DOUT_TEMPR71[9] , \A_DOUT_TEMPR71[8] , 
        \A_DOUT_TEMPR71[7] , \A_DOUT_TEMPR71[6] , \A_DOUT_TEMPR71[5] })
        , .B_DOUT({nc1905, nc1906, nc1907, nc1908, nc1909, nc1910, 
        nc1911, nc1912, nc1913, nc1914, nc1915, nc1916, nc1917, nc1918, 
        nc1919, \B_DOUT_TEMPR71[9] , \B_DOUT_TEMPR71[8] , 
        \B_DOUT_TEMPR71[7] , \B_DOUT_TEMPR71[6] , \B_DOUT_TEMPR71[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[71][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_209 (.A(\B_DOUT_TEMPR28[0] ), .B(\B_DOUT_TEMPR29[0] ), .C(
        \B_DOUT_TEMPR30[0] ), .D(\B_DOUT_TEMPR31[0] ), .Y(OR4_209_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%92%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R92C1 (
        .A_DOUT({nc1920, nc1921, nc1922, nc1923, nc1924, nc1925, 
        nc1926, nc1927, nc1928, nc1929, nc1930, nc1931, nc1932, nc1933, 
        nc1934, \A_DOUT_TEMPR92[9] , \A_DOUT_TEMPR92[8] , 
        \A_DOUT_TEMPR92[7] , \A_DOUT_TEMPR92[6] , \A_DOUT_TEMPR92[5] })
        , .B_DOUT({nc1935, nc1936, nc1937, nc1938, nc1939, nc1940, 
        nc1941, nc1942, nc1943, nc1944, nc1945, nc1946, nc1947, nc1948, 
        nc1949, \B_DOUT_TEMPR92[9] , \B_DOUT_TEMPR92[8] , 
        \B_DOUT_TEMPR92[7] , \B_DOUT_TEMPR92[6] , \B_DOUT_TEMPR92[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[92][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1323 (.A(\A_DOUT_TEMPR20[21] ), .B(\A_DOUT_TEMPR21[21] ), 
        .C(\A_DOUT_TEMPR22[21] ), .D(\A_DOUT_TEMPR23[21] ), .Y(
        OR4_1323_Y));
    OR4 OR4_2042 (.A(\A_DOUT_TEMPR48[0] ), .B(\A_DOUT_TEMPR49[0] ), .C(
        \A_DOUT_TEMPR50[0] ), .D(\A_DOUT_TEMPR51[0] ), .Y(OR4_2042_Y));
    OR4 OR4_2402 (.A(\B_DOUT_TEMPR99[7] ), .B(\B_DOUT_TEMPR100[7] ), 
        .C(\B_DOUT_TEMPR101[7] ), .D(\B_DOUT_TEMPR102[7] ), .Y(
        OR4_2402_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%102%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R102C7 (
        .A_DOUT({nc1950, nc1951, nc1952, nc1953, nc1954, nc1955, 
        nc1956, nc1957, nc1958, nc1959, nc1960, nc1961, nc1962, nc1963, 
        nc1964, \A_DOUT_TEMPR102[39] , \A_DOUT_TEMPR102[38] , 
        \A_DOUT_TEMPR102[37] , \A_DOUT_TEMPR102[36] , 
        \A_DOUT_TEMPR102[35] }), .B_DOUT({nc1965, nc1966, nc1967, 
        nc1968, nc1969, nc1970, nc1971, nc1972, nc1973, nc1974, nc1975, 
        nc1976, nc1977, nc1978, nc1979, \B_DOUT_TEMPR102[39] , 
        \B_DOUT_TEMPR102[38] , \B_DOUT_TEMPR102[37] , 
        \B_DOUT_TEMPR102[36] , \B_DOUT_TEMPR102[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[102][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h40) )  CFG3_20 (.A(B_ADDR[16]), .B(B_ADDR[15]), 
        .C(B_ADDR[14]), .Y(CFG3_20_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%84%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R84C2 (
        .A_DOUT({nc1980, nc1981, nc1982, nc1983, nc1984, nc1985, 
        nc1986, nc1987, nc1988, nc1989, nc1990, nc1991, nc1992, nc1993, 
        nc1994, \A_DOUT_TEMPR84[14] , \A_DOUT_TEMPR84[13] , 
        \A_DOUT_TEMPR84[12] , \A_DOUT_TEMPR84[11] , 
        \A_DOUT_TEMPR84[10] }), .B_DOUT({nc1995, nc1996, nc1997, 
        nc1998, nc1999, nc2000, nc2001, nc2002, nc2003, nc2004, nc2005, 
        nc2006, nc2007, nc2008, nc2009, \B_DOUT_TEMPR84[14] , 
        \B_DOUT_TEMPR84[13] , \B_DOUT_TEMPR84[12] , 
        \B_DOUT_TEMPR84[11] , \B_DOUT_TEMPR84[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[84][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[17]  (.A(OR4_440_Y), .B(OR4_2199_Y), .C(OR4_1231_Y)
        , .D(OR4_2378_Y), .Y(A_DOUT[17]));
    OR4 OR4_703 (.A(\A_DOUT_TEMPR95[6] ), .B(\A_DOUT_TEMPR96[6] ), .C(
        \A_DOUT_TEMPR97[6] ), .D(\A_DOUT_TEMPR98[6] ), .Y(OR4_703_Y));
    OR4 OR4_488 (.A(\B_DOUT_TEMPR12[13] ), .B(\B_DOUT_TEMPR13[13] ), 
        .C(\B_DOUT_TEMPR14[13] ), .D(\B_DOUT_TEMPR15[13] ), .Y(
        OR4_488_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%43%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R43C2 (
        .A_DOUT({nc2010, nc2011, nc2012, nc2013, nc2014, nc2015, 
        nc2016, nc2017, nc2018, nc2019, nc2020, nc2021, nc2022, nc2023, 
        nc2024, \A_DOUT_TEMPR43[14] , \A_DOUT_TEMPR43[13] , 
        \A_DOUT_TEMPR43[12] , \A_DOUT_TEMPR43[11] , 
        \A_DOUT_TEMPR43[10] }), .B_DOUT({nc2025, nc2026, nc2027, 
        nc2028, nc2029, nc2030, nc2031, nc2032, nc2033, nc2034, nc2035, 
        nc2036, nc2037, nc2038, nc2039, \B_DOUT_TEMPR43[14] , 
        \B_DOUT_TEMPR43[13] , \B_DOUT_TEMPR43[12] , 
        \B_DOUT_TEMPR43[11] , \B_DOUT_TEMPR43[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[43][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2408 (.A(\B_DOUT_TEMPR4[11] ), .B(\B_DOUT_TEMPR5[11] ), .C(
        \B_DOUT_TEMPR6[11] ), .D(\B_DOUT_TEMPR7[11] ), .Y(OR4_2408_Y));
    OR4 OR4_1365 (.A(OR4_104_Y), .B(OR4_1599_Y), .C(OR4_2166_Y), .D(
        OR4_1999_Y), .Y(OR4_1365_Y));
    OR4 OR4_584 (.A(\B_DOUT_TEMPR4[14] ), .B(\B_DOUT_TEMPR5[14] ), .C(
        \B_DOUT_TEMPR6[14] ), .D(\B_DOUT_TEMPR7[14] ), .Y(OR4_584_Y));
    OR4 OR4_27 (.A(\A_DOUT_TEMPR28[23] ), .B(\A_DOUT_TEMPR29[23] ), .C(
        \A_DOUT_TEMPR30[23] ), .D(\A_DOUT_TEMPR31[23] ), .Y(OR4_27_Y));
    OR4 OR4_731 (.A(\B_DOUT_TEMPR115[8] ), .B(\B_DOUT_TEMPR116[8] ), 
        .C(\B_DOUT_TEMPR117[8] ), .D(\B_DOUT_TEMPR118[8] ), .Y(
        OR4_731_Y));
    OR4 OR4_116 (.A(OR4_133_Y), .B(OR4_531_Y), .C(OR4_1291_Y), .D(
        OR4_2092_Y), .Y(OR4_116_Y));
    OR4 OR4_177 (.A(\B_DOUT_TEMPR95[37] ), .B(\B_DOUT_TEMPR96[37] ), 
        .C(\B_DOUT_TEMPR97[37] ), .D(\B_DOUT_TEMPR98[37] ), .Y(
        OR4_177_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%2%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R2C4 (
        .A_DOUT({nc2040, nc2041, nc2042, nc2043, nc2044, nc2045, 
        nc2046, nc2047, nc2048, nc2049, nc2050, nc2051, nc2052, nc2053, 
        nc2054, \A_DOUT_TEMPR2[24] , \A_DOUT_TEMPR2[23] , 
        \A_DOUT_TEMPR2[22] , \A_DOUT_TEMPR2[21] , \A_DOUT_TEMPR2[20] })
        , .B_DOUT({nc2055, nc2056, nc2057, nc2058, nc2059, nc2060, 
        nc2061, nc2062, nc2063, nc2064, nc2065, nc2066, nc2067, nc2068, 
        nc2069, \B_DOUT_TEMPR2[24] , \B_DOUT_TEMPR2[23] , 
        \B_DOUT_TEMPR2[22] , \B_DOUT_TEMPR2[21] , \B_DOUT_TEMPR2[20] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[2][4] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[24], A_DIN[23], A_DIN[22], 
        A_DIN[21], A_DIN[20]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%55%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R55C2 (
        .A_DOUT({nc2070, nc2071, nc2072, nc2073, nc2074, nc2075, 
        nc2076, nc2077, nc2078, nc2079, nc2080, nc2081, nc2082, nc2083, 
        nc2084, \A_DOUT_TEMPR55[14] , \A_DOUT_TEMPR55[13] , 
        \A_DOUT_TEMPR55[12] , \A_DOUT_TEMPR55[11] , 
        \A_DOUT_TEMPR55[10] }), .B_DOUT({nc2085, nc2086, nc2087, 
        nc2088, nc2089, nc2090, nc2091, nc2092, nc2093, nc2094, nc2095, 
        nc2096, nc2097, nc2098, nc2099, \B_DOUT_TEMPR55[14] , 
        \B_DOUT_TEMPR55[13] , \B_DOUT_TEMPR55[12] , 
        \B_DOUT_TEMPR55[11] , \B_DOUT_TEMPR55[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[55][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1445 (.A(OR4_1029_Y), .B(OR4_1849_Y), .C(OR4_285_Y), .D(
        OR4_1854_Y), .Y(OR4_1445_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%1%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R1C1 (
        .A_DOUT({nc2100, nc2101, nc2102, nc2103, nc2104, nc2105, 
        nc2106, nc2107, nc2108, nc2109, nc2110, nc2111, nc2112, nc2113, 
        nc2114, \A_DOUT_TEMPR1[9] , \A_DOUT_TEMPR1[8] , 
        \A_DOUT_TEMPR1[7] , \A_DOUT_TEMPR1[6] , \A_DOUT_TEMPR1[5] }), 
        .B_DOUT({nc2115, nc2116, nc2117, nc2118, nc2119, nc2120, 
        nc2121, nc2122, nc2123, nc2124, nc2125, nc2126, nc2127, nc2128, 
        nc2129, \B_DOUT_TEMPR1[9] , \B_DOUT_TEMPR1[8] , 
        \B_DOUT_TEMPR1[7] , \B_DOUT_TEMPR1[6] , \B_DOUT_TEMPR1[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[1][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[0] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[0] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%14%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R14C3 (
        .A_DOUT({nc2130, nc2131, nc2132, nc2133, nc2134, nc2135, 
        nc2136, nc2137, nc2138, nc2139, nc2140, nc2141, nc2142, nc2143, 
        nc2144, \A_DOUT_TEMPR14[19] , \A_DOUT_TEMPR14[18] , 
        \A_DOUT_TEMPR14[17] , \A_DOUT_TEMPR14[16] , 
        \A_DOUT_TEMPR14[15] }), .B_DOUT({nc2145, nc2146, nc2147, 
        nc2148, nc2149, nc2150, nc2151, nc2152, nc2153, nc2154, nc2155, 
        nc2156, nc2157, nc2158, nc2159, \B_DOUT_TEMPR14[19] , 
        \B_DOUT_TEMPR14[18] , \B_DOUT_TEMPR14[17] , 
        \B_DOUT_TEMPR14[16] , \B_DOUT_TEMPR14[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[14][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_208 (.A(\A_DOUT_TEMPR107[30] ), .B(\A_DOUT_TEMPR108[30] ), 
        .C(\A_DOUT_TEMPR109[30] ), .D(\A_DOUT_TEMPR110[30] ), .Y(
        OR4_208_Y));
    OR4 OR4_1502 (.A(\A_DOUT_TEMPR68[28] ), .B(\A_DOUT_TEMPR69[28] ), 
        .C(\A_DOUT_TEMPR70[28] ), .D(\A_DOUT_TEMPR71[28] ), .Y(
        OR4_1502_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%83%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R83C7 (
        .A_DOUT({nc2160, nc2161, nc2162, nc2163, nc2164, nc2165, 
        nc2166, nc2167, nc2168, nc2169, nc2170, nc2171, nc2172, nc2173, 
        nc2174, \A_DOUT_TEMPR83[39] , \A_DOUT_TEMPR83[38] , 
        \A_DOUT_TEMPR83[37] , \A_DOUT_TEMPR83[36] , 
        \A_DOUT_TEMPR83[35] }), .B_DOUT({nc2175, nc2176, nc2177, 
        nc2178, nc2179, nc2180, nc2181, nc2182, nc2183, nc2184, nc2185, 
        nc2186, nc2187, nc2188, nc2189, \B_DOUT_TEMPR83[39] , 
        \B_DOUT_TEMPR83[38] , \B_DOUT_TEMPR83[37] , 
        \B_DOUT_TEMPR83[36] , \B_DOUT_TEMPR83[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[83][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2500 (.A(\B_DOUT_TEMPR44[12] ), .B(\B_DOUT_TEMPR45[12] ), 
        .C(\B_DOUT_TEMPR46[12] ), .D(\B_DOUT_TEMPR47[12] ), .Y(
        OR4_2500_Y));
    OR2 OR2_63 (.A(\B_DOUT_TEMPR72[29] ), .B(\B_DOUT_TEMPR73[29] ), .Y(
        OR2_63_Y));
    OR4 OR4_2973 (.A(\B_DOUT_TEMPR44[30] ), .B(\B_DOUT_TEMPR45[30] ), 
        .C(\B_DOUT_TEMPR46[30] ), .D(\B_DOUT_TEMPR47[30] ), .Y(
        OR4_2973_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENA[8]  (.A(A_WBYTE_EN[4]), .B(
        A_WEN), .Y(\WBYTEENA[8] ));
    OR4 OR4_1594 (.A(OR4_1281_Y), .B(OR4_1570_Y), .C(OR4_1224_Y), .D(
        OR4_1582_Y), .Y(OR4_1594_Y));
    OR4 OR4_832 (.A(\B_DOUT_TEMPR107[23] ), .B(\B_DOUT_TEMPR108[23] ), 
        .C(\B_DOUT_TEMPR109[23] ), .D(\B_DOUT_TEMPR110[23] ), .Y(
        OR4_832_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%62%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R62C6 (
        .A_DOUT({nc2190, nc2191, nc2192, nc2193, nc2194, nc2195, 
        nc2196, nc2197, nc2198, nc2199, nc2200, nc2201, nc2202, nc2203, 
        nc2204, \A_DOUT_TEMPR62[34] , \A_DOUT_TEMPR62[33] , 
        \A_DOUT_TEMPR62[32] , \A_DOUT_TEMPR62[31] , 
        \A_DOUT_TEMPR62[30] }), .B_DOUT({nc2205, nc2206, nc2207, 
        nc2208, nc2209, nc2210, nc2211, nc2212, nc2213, nc2214, nc2215, 
        nc2216, nc2217, nc2218, nc2219, \B_DOUT_TEMPR62[34] , 
        \B_DOUT_TEMPR62[33] , \B_DOUT_TEMPR62[32] , 
        \B_DOUT_TEMPR62[31] , \B_DOUT_TEMPR62[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[62][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1781 (.A(OR4_2020_Y), .B(OR4_402_Y), .C(OR2_77_Y), .D(
        \A_DOUT_TEMPR74[2] ), .Y(OR4_1781_Y));
    OR2 OR2_13 (.A(\A_DOUT_TEMPR72[3] ), .B(\A_DOUT_TEMPR73[3] ), .Y(
        OR2_13_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%49%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R49C4 (
        .A_DOUT({nc2220, nc2221, nc2222, nc2223, nc2224, nc2225, 
        nc2226, nc2227, nc2228, nc2229, nc2230, nc2231, nc2232, nc2233, 
        nc2234, \A_DOUT_TEMPR49[24] , \A_DOUT_TEMPR49[23] , 
        \A_DOUT_TEMPR49[22] , \A_DOUT_TEMPR49[21] , 
        \A_DOUT_TEMPR49[20] }), .B_DOUT({nc2235, nc2236, nc2237, 
        nc2238, nc2239, nc2240, nc2241, nc2242, nc2243, nc2244, nc2245, 
        nc2246, nc2247, nc2248, nc2249, \B_DOUT_TEMPR49[24] , 
        \B_DOUT_TEMPR49[23] , \B_DOUT_TEMPR49[22] , 
        \B_DOUT_TEMPR49[21] , \B_DOUT_TEMPR49[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[49][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1517 (.A(\B_DOUT_TEMPR48[24] ), .B(\B_DOUT_TEMPR49[24] ), 
        .C(\B_DOUT_TEMPR50[24] ), .D(\B_DOUT_TEMPR51[24] ), .Y(
        OR4_1517_Y));
    OR4 OR4_2819 (.A(OR4_1065_Y), .B(OR4_1356_Y), .C(OR4_2962_Y), .D(
        OR4_826_Y), .Y(OR4_2819_Y));
    OR4 OR4_1746 (.A(\B_DOUT_TEMPR107[11] ), .B(\B_DOUT_TEMPR108[11] ), 
        .C(\B_DOUT_TEMPR109[11] ), .D(\B_DOUT_TEMPR110[11] ), .Y(
        OR4_1746_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%69%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R69C0 (
        .A_DOUT({nc2250, nc2251, nc2252, nc2253, nc2254, nc2255, 
        nc2256, nc2257, nc2258, nc2259, nc2260, nc2261, nc2262, nc2263, 
        nc2264, \A_DOUT_TEMPR69[4] , \A_DOUT_TEMPR69[3] , 
        \A_DOUT_TEMPR69[2] , \A_DOUT_TEMPR69[1] , \A_DOUT_TEMPR69[0] })
        , .B_DOUT({nc2265, nc2266, nc2267, nc2268, nc2269, nc2270, 
        nc2271, nc2272, nc2273, nc2274, nc2275, nc2276, nc2277, nc2278, 
        nc2279, \B_DOUT_TEMPR69[4] , \B_DOUT_TEMPR69[3] , 
        \B_DOUT_TEMPR69[2] , \B_DOUT_TEMPR69[1] , \B_DOUT_TEMPR69[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[69][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_513 (.A(\B_DOUT_TEMPR99[4] ), .B(\B_DOUT_TEMPR100[4] ), .C(
        \B_DOUT_TEMPR101[4] ), .D(\B_DOUT_TEMPR102[4] ), .Y(OR4_513_Y));
    OR4 OR4_20 (.A(\B_DOUT_TEMPR52[3] ), .B(\B_DOUT_TEMPR53[3] ), .C(
        \B_DOUT_TEMPR54[3] ), .D(\B_DOUT_TEMPR55[3] ), .Y(OR4_20_Y));
    OR4 OR4_2371 (.A(\A_DOUT_TEMPR83[20] ), .B(\A_DOUT_TEMPR84[20] ), 
        .C(\A_DOUT_TEMPR85[20] ), .D(\A_DOUT_TEMPR86[20] ), .Y(
        OR4_2371_Y));
    OR4 OR4_1953 (.A(\B_DOUT_TEMPR79[19] ), .B(\B_DOUT_TEMPR80[19] ), 
        .C(\B_DOUT_TEMPR81[19] ), .D(\B_DOUT_TEMPR82[19] ), .Y(
        OR4_1953_Y));
    OR4 OR4_2111 (.A(\B_DOUT_TEMPR68[17] ), .B(\B_DOUT_TEMPR69[17] ), 
        .C(\B_DOUT_TEMPR70[17] ), .D(\B_DOUT_TEMPR71[17] ), .Y(
        OR4_2111_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%65%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R65C6 (
        .A_DOUT({nc2280, nc2281, nc2282, nc2283, nc2284, nc2285, 
        nc2286, nc2287, nc2288, nc2289, nc2290, nc2291, nc2292, nc2293, 
        nc2294, \A_DOUT_TEMPR65[34] , \A_DOUT_TEMPR65[33] , 
        \A_DOUT_TEMPR65[32] , \A_DOUT_TEMPR65[31] , 
        \A_DOUT_TEMPR65[30] }), .B_DOUT({nc2295, nc2296, nc2297, 
        nc2298, nc2299, nc2300, nc2301, nc2302, nc2303, nc2304, nc2305, 
        nc2306, nc2307, nc2308, nc2309, \B_DOUT_TEMPR65[34] , 
        \B_DOUT_TEMPR65[33] , \B_DOUT_TEMPR65[32] , 
        \B_DOUT_TEMPR65[31] , \B_DOUT_TEMPR65[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[65][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_107 (.A(\A_DOUT_TEMPR0[24] ), .B(\A_DOUT_TEMPR1[24] ), .C(
        \A_DOUT_TEMPR2[24] ), .D(\A_DOUT_TEMPR3[24] ), .Y(OR4_107_Y));
    OR4 OR4_15 (.A(\A_DOUT_TEMPR16[26] ), .B(\A_DOUT_TEMPR17[26] ), .C(
        \A_DOUT_TEMPR18[26] ), .D(\A_DOUT_TEMPR19[26] ), .Y(OR4_15_Y));
    OR4 OR4_759 (.A(\B_DOUT_TEMPR60[26] ), .B(\B_DOUT_TEMPR61[26] ), 
        .C(\B_DOUT_TEMPR62[26] ), .D(\B_DOUT_TEMPR63[26] ), .Y(
        OR4_759_Y));
    OR4 OR4_2871 (.A(\A_DOUT_TEMPR48[33] ), .B(\A_DOUT_TEMPR49[33] ), 
        .C(\A_DOUT_TEMPR50[33] ), .D(\A_DOUT_TEMPR51[33] ), .Y(
        OR4_2871_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%21%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R21C5 (
        .A_DOUT({nc2310, nc2311, nc2312, nc2313, nc2314, nc2315, 
        nc2316, nc2317, nc2318, nc2319, nc2320, nc2321, nc2322, nc2323, 
        nc2324, \A_DOUT_TEMPR21[29] , \A_DOUT_TEMPR21[28] , 
        \A_DOUT_TEMPR21[27] , \A_DOUT_TEMPR21[26] , 
        \A_DOUT_TEMPR21[25] }), .B_DOUT({nc2325, nc2326, nc2327, 
        nc2328, nc2329, nc2330, nc2331, nc2332, nc2333, nc2334, nc2335, 
        nc2336, nc2337, nc2338, nc2339, \B_DOUT_TEMPR21[29] , 
        \B_DOUT_TEMPR21[28] , \B_DOUT_TEMPR21[27] , 
        \B_DOUT_TEMPR21[26] , \B_DOUT_TEMPR21[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[21][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[34]  (.A(OR4_2940_Y), .B(OR4_1526_Y), .C(
        OR4_1696_Y), .D(OR4_2970_Y), .Y(A_DOUT[34]));
    OR4 OR4_589 (.A(\A_DOUT_TEMPR60[37] ), .B(\A_DOUT_TEMPR61[37] ), 
        .C(\A_DOUT_TEMPR62[37] ), .D(\A_DOUT_TEMPR63[37] ), .Y(
        OR4_589_Y));
    OR4 OR4_1291 (.A(\A_DOUT_TEMPR24[28] ), .B(\A_DOUT_TEMPR25[28] ), 
        .C(\A_DOUT_TEMPR26[28] ), .D(\A_DOUT_TEMPR27[28] ), .Y(
        OR4_1291_Y));
    OR4 OR4_2015 (.A(OR4_2044_Y), .B(OR4_1857_Y), .C(OR4_1795_Y), .D(
        OR4_74_Y), .Y(OR4_2015_Y));
    OR4 OR4_655 (.A(\A_DOUT_TEMPR36[2] ), .B(\A_DOUT_TEMPR37[2] ), .C(
        \A_DOUT_TEMPR38[2] ), .D(\A_DOUT_TEMPR39[2] ), .Y(OR4_655_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%108%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R108C4 (
        .A_DOUT({nc2340, nc2341, nc2342, nc2343, nc2344, nc2345, 
        nc2346, nc2347, nc2348, nc2349, nc2350, nc2351, nc2352, nc2353, 
        nc2354, \A_DOUT_TEMPR108[24] , \A_DOUT_TEMPR108[23] , 
        \A_DOUT_TEMPR108[22] , \A_DOUT_TEMPR108[21] , 
        \A_DOUT_TEMPR108[20] }), .B_DOUT({nc2355, nc2356, nc2357, 
        nc2358, nc2359, nc2360, nc2361, nc2362, nc2363, nc2364, nc2365, 
        nc2366, nc2367, nc2368, nc2369, \B_DOUT_TEMPR108[24] , 
        \B_DOUT_TEMPR108[23] , \B_DOUT_TEMPR108[22] , 
        \B_DOUT_TEMPR108[21] , \B_DOUT_TEMPR108[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[108][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2557 (.A(\A_DOUT_TEMPR36[38] ), .B(\A_DOUT_TEMPR37[38] ), 
        .C(\A_DOUT_TEMPR38[38] ), .D(\A_DOUT_TEMPR39[38] ), .Y(
        OR4_2557_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%35%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R35C2 (
        .A_DOUT({nc2370, nc2371, nc2372, nc2373, nc2374, nc2375, 
        nc2376, nc2377, nc2378, nc2379, nc2380, nc2381, nc2382, nc2383, 
        nc2384, \A_DOUT_TEMPR35[14] , \A_DOUT_TEMPR35[13] , 
        \A_DOUT_TEMPR35[12] , \A_DOUT_TEMPR35[11] , 
        \A_DOUT_TEMPR35[10] }), .B_DOUT({nc2385, nc2386, nc2387, 
        nc2388, nc2389, nc2390, nc2391, nc2392, nc2393, nc2394, nc2395, 
        nc2396, nc2397, nc2398, nc2399, \B_DOUT_TEMPR35[14] , 
        \B_DOUT_TEMPR35[13] , \B_DOUT_TEMPR35[12] , 
        \B_DOUT_TEMPR35[11] , \B_DOUT_TEMPR35[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[35][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2905 (.A(\B_DOUT_TEMPR64[33] ), .B(\B_DOUT_TEMPR65[33] ), 
        .C(\B_DOUT_TEMPR66[33] ), .D(\B_DOUT_TEMPR67[33] ), .Y(
        OR4_2905_Y));
    OR4 OR4_259 (.A(\B_DOUT_TEMPR32[20] ), .B(\B_DOUT_TEMPR33[20] ), 
        .C(\B_DOUT_TEMPR34[20] ), .D(\B_DOUT_TEMPR35[20] ), .Y(
        OR4_259_Y));
    OR4 OR4_1351 (.A(\A_DOUT_TEMPR56[6] ), .B(\A_DOUT_TEMPR57[6] ), .C(
        \A_DOUT_TEMPR58[6] ), .D(\A_DOUT_TEMPR59[6] ), .Y(OR4_1351_Y));
    OR4 OR4_1000 (.A(OR4_3029_Y), .B(OR4_2177_Y), .C(OR4_1195_Y), .D(
        OR4_1465_Y), .Y(OR4_1000_Y));
    OR4 OR4_2721 (.A(\A_DOUT_TEMPR68[19] ), .B(\A_DOUT_TEMPR69[19] ), 
        .C(\A_DOUT_TEMPR70[19] ), .D(\A_DOUT_TEMPR71[19] ), .Y(
        OR4_2721_Y));
    OR4 OR4_1483 (.A(\B_DOUT_TEMPR115[32] ), .B(\B_DOUT_TEMPR116[32] ), 
        .C(\B_DOUT_TEMPR117[32] ), .D(\B_DOUT_TEMPR118[32] ), .Y(
        OR4_1483_Y));
    OR4 OR4_1851 (.A(\B_DOUT_TEMPR111[15] ), .B(\B_DOUT_TEMPR112[15] ), 
        .C(\B_DOUT_TEMPR113[15] ), .D(\B_DOUT_TEMPR114[15] ), .Y(
        OR4_1851_Y));
    OR4 OR4_2609 (.A(OR4_346_Y), .B(OR4_2403_Y), .C(OR4_2627_Y), .D(
        OR4_2417_Y), .Y(OR4_2609_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%83%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R83C0 (
        .A_DOUT({nc2400, nc2401, nc2402, nc2403, nc2404, nc2405, 
        nc2406, nc2407, nc2408, nc2409, nc2410, nc2411, nc2412, nc2413, 
        nc2414, \A_DOUT_TEMPR83[4] , \A_DOUT_TEMPR83[3] , 
        \A_DOUT_TEMPR83[2] , \A_DOUT_TEMPR83[1] , \A_DOUT_TEMPR83[0] })
        , .B_DOUT({nc2415, nc2416, nc2417, nc2418, nc2419, nc2420, 
        nc2421, nc2422, nc2423, nc2424, nc2425, nc2426, nc2427, nc2428, 
        nc2429, \B_DOUT_TEMPR83[4] , \B_DOUT_TEMPR83[3] , 
        \B_DOUT_TEMPR83[2] , \B_DOUT_TEMPR83[1] , \B_DOUT_TEMPR83[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[83][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_753 (.A(OR4_1762_Y), .B(OR4_56_Y), .C(OR4_2758_Y), .D(
        OR4_739_Y), .Y(OR4_753_Y));
    OR4 OR4_276 (.A(OR4_459_Y), .B(OR4_2497_Y), .C(OR4_966_Y), .D(
        OR4_2500_Y), .Y(OR4_276_Y));
    OR4 OR4_2817 (.A(\A_DOUT_TEMPR56[3] ), .B(\A_DOUT_TEMPR57[3] ), .C(
        \A_DOUT_TEMPR58[3] ), .D(\A_DOUT_TEMPR59[3] ), .Y(OR4_2817_Y));
    OR4 OR4_2139 (.A(\A_DOUT_TEMPR87[34] ), .B(\A_DOUT_TEMPR88[34] ), 
        .C(\A_DOUT_TEMPR89[34] ), .D(\A_DOUT_TEMPR90[34] ), .Y(
        OR4_2139_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%113%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R113C7 (
        .A_DOUT({nc2430, nc2431, nc2432, nc2433, nc2434, nc2435, 
        nc2436, nc2437, nc2438, nc2439, nc2440, nc2441, nc2442, nc2443, 
        nc2444, \A_DOUT_TEMPR113[39] , \A_DOUT_TEMPR113[38] , 
        \A_DOUT_TEMPR113[37] , \A_DOUT_TEMPR113[36] , 
        \A_DOUT_TEMPR113[35] }), .B_DOUT({nc2445, nc2446, nc2447, 
        nc2448, nc2449, nc2450, nc2451, nc2452, nc2453, nc2454, nc2455, 
        nc2456, nc2457, nc2458, nc2459, \B_DOUT_TEMPR113[39] , 
        \B_DOUT_TEMPR113[38] , \B_DOUT_TEMPR113[37] , 
        \B_DOUT_TEMPR113[36] , \B_DOUT_TEMPR113[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[113][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1218 (.A(\A_DOUT_TEMPR83[2] ), .B(\A_DOUT_TEMPR84[2] ), .C(
        \A_DOUT_TEMPR85[2] ), .D(\A_DOUT_TEMPR86[2] ), .Y(OR4_1218_Y));
    OR4 OR4_1139 (.A(OR4_1780_Y), .B(OR4_1590_Y), .C(OR4_2457_Y), .D(
        OR4_617_Y), .Y(OR4_1139_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%3%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R3C2 (
        .A_DOUT({nc2460, nc2461, nc2462, nc2463, nc2464, nc2465, 
        nc2466, nc2467, nc2468, nc2469, nc2470, nc2471, nc2472, nc2473, 
        nc2474, \A_DOUT_TEMPR3[14] , \A_DOUT_TEMPR3[13] , 
        \A_DOUT_TEMPR3[12] , \A_DOUT_TEMPR3[11] , \A_DOUT_TEMPR3[10] })
        , .B_DOUT({nc2475, nc2476, nc2477, nc2478, nc2479, nc2480, 
        nc2481, nc2482, nc2483, nc2484, nc2485, nc2486, nc2487, nc2488, 
        nc2489, \B_DOUT_TEMPR3[14] , \B_DOUT_TEMPR3[13] , 
        \B_DOUT_TEMPR3[12] , \B_DOUT_TEMPR3[11] , \B_DOUT_TEMPR3[10] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[3][2] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[14], A_DIN[13], A_DIN[12], 
        A_DIN[11], A_DIN[10]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_258 (.A(OR4_1205_Y), .B(OR4_2694_Y), .C(OR4_215_Y), .D(
        OR4_44_Y), .Y(OR4_258_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%87%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R87C7 (
        .A_DOUT({nc2490, nc2491, nc2492, nc2493, nc2494, nc2495, 
        nc2496, nc2497, nc2498, nc2499, nc2500, nc2501, nc2502, nc2503, 
        nc2504, \A_DOUT_TEMPR87[39] , \A_DOUT_TEMPR87[38] , 
        \A_DOUT_TEMPR87[37] , \A_DOUT_TEMPR87[36] , 
        \A_DOUT_TEMPR87[35] }), .B_DOUT({nc2505, nc2506, nc2507, 
        nc2508, nc2509, nc2510, nc2511, nc2512, nc2513, nc2514, nc2515, 
        nc2516, nc2517, nc2518, nc2519, \B_DOUT_TEMPR87[39] , 
        \B_DOUT_TEMPR87[38] , \B_DOUT_TEMPR87[37] , 
        \B_DOUT_TEMPR87[36] , \B_DOUT_TEMPR87[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[87][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%52%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R52C5 (
        .A_DOUT({nc2520, nc2521, nc2522, nc2523, nc2524, nc2525, 
        nc2526, nc2527, nc2528, nc2529, nc2530, nc2531, nc2532, nc2533, 
        nc2534, \A_DOUT_TEMPR52[29] , \A_DOUT_TEMPR52[28] , 
        \A_DOUT_TEMPR52[27] , \A_DOUT_TEMPR52[26] , 
        \A_DOUT_TEMPR52[25] }), .B_DOUT({nc2535, nc2536, nc2537, 
        nc2538, nc2539, nc2540, nc2541, nc2542, nc2543, nc2544, nc2545, 
        nc2546, nc2547, nc2548, nc2549, \B_DOUT_TEMPR52[29] , 
        \B_DOUT_TEMPR52[28] , \B_DOUT_TEMPR52[27] , 
        \B_DOUT_TEMPR52[26] , \B_DOUT_TEMPR52[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[52][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%114%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R114C7 (
        .A_DOUT({nc2550, nc2551, nc2552, nc2553, nc2554, nc2555, 
        nc2556, nc2557, nc2558, nc2559, nc2560, nc2561, nc2562, nc2563, 
        nc2564, \A_DOUT_TEMPR114[39] , \A_DOUT_TEMPR114[38] , 
        \A_DOUT_TEMPR114[37] , \A_DOUT_TEMPR114[36] , 
        \A_DOUT_TEMPR114[35] }), .B_DOUT({nc2565, nc2566, nc2567, 
        nc2568, nc2569, nc2570, nc2571, nc2572, nc2573, nc2574, nc2575, 
        nc2576, nc2577, nc2578, nc2579, \B_DOUT_TEMPR114[39] , 
        \B_DOUT_TEMPR114[38] , \B_DOUT_TEMPR114[37] , 
        \B_DOUT_TEMPR114[36] , \B_DOUT_TEMPR114[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[114][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2348 (.A(\A_DOUT_TEMPR12[39] ), .B(\A_DOUT_TEMPR13[39] ), 
        .C(\A_DOUT_TEMPR14[39] ), .D(\A_DOUT_TEMPR15[39] ), .Y(
        OR4_2348_Y));
    OR4 \OR4_B_DOUT[31]  (.A(OR4_1137_Y), .B(OR4_675_Y), .C(OR4_2021_Y)
        , .D(OR4_1010_Y), .Y(B_DOUT[31]));
    OR4 OR4_737 (.A(OR4_124_Y), .B(OR4_1335_Y), .C(OR2_56_Y), .D(
        \B_DOUT_TEMPR74[18] ), .Y(OR4_737_Y));
    OR4 \OR4_A_DOUT[2]  (.A(OR4_2713_Y), .B(OR4_319_Y), .C(OR4_349_Y), 
        .D(OR4_754_Y), .Y(A_DOUT[2]));
    OR4 OR4_333 (.A(\B_DOUT_TEMPR40[29] ), .B(\B_DOUT_TEMPR41[29] ), 
        .C(\B_DOUT_TEMPR42[29] ), .D(\B_DOUT_TEMPR43[29] ), .Y(
        OR4_333_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%52%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R52C1 (
        .A_DOUT({nc2580, nc2581, nc2582, nc2583, nc2584, nc2585, 
        nc2586, nc2587, nc2588, nc2589, nc2590, nc2591, nc2592, nc2593, 
        nc2594, \A_DOUT_TEMPR52[9] , \A_DOUT_TEMPR52[8] , 
        \A_DOUT_TEMPR52[7] , \A_DOUT_TEMPR52[6] , \A_DOUT_TEMPR52[5] })
        , .B_DOUT({nc2595, nc2596, nc2597, nc2598, nc2599, nc2600, 
        nc2601, nc2602, nc2603, nc2604, nc2605, nc2606, nc2607, nc2608, 
        nc2609, \B_DOUT_TEMPR52[9] , \B_DOUT_TEMPR52[8] , 
        \B_DOUT_TEMPR52[7] , \B_DOUT_TEMPR52[6] , \B_DOUT_TEMPR52[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[52][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2423 (.A(\B_DOUT_TEMPR83[39] ), .B(\B_DOUT_TEMPR84[39] ), 
        .C(\B_DOUT_TEMPR85[39] ), .D(\B_DOUT_TEMPR86[39] ), .Y(
        OR4_2423_Y));
    OR4 OR4_166 (.A(\B_DOUT_TEMPR52[9] ), .B(\B_DOUT_TEMPR53[9] ), .C(
        \B_DOUT_TEMPR54[9] ), .D(\B_DOUT_TEMPR55[9] ), .Y(OR4_166_Y));
    OR4 OR4_738 (.A(OR4_92_Y), .B(OR4_943_Y), .C(OR2_79_Y), .D(
        \B_DOUT_TEMPR74[20] ), .Y(OR4_738_Y));
    OR4 OR4_1406 (.A(\B_DOUT_TEMPR40[8] ), .B(\B_DOUT_TEMPR41[8] ), .C(
        \B_DOUT_TEMPR42[8] ), .D(\B_DOUT_TEMPR43[8] ), .Y(OR4_1406_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%6%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R6C1 (
        .A_DOUT({nc2610, nc2611, nc2612, nc2613, nc2614, nc2615, 
        nc2616, nc2617, nc2618, nc2619, nc2620, nc2621, nc2622, nc2623, 
        nc2624, \A_DOUT_TEMPR6[9] , \A_DOUT_TEMPR6[8] , 
        \A_DOUT_TEMPR6[7] , \A_DOUT_TEMPR6[6] , \A_DOUT_TEMPR6[5] }), 
        .B_DOUT({nc2625, nc2626, nc2627, nc2628, nc2629, nc2630, 
        nc2631, nc2632, nc2633, nc2634, nc2635, nc2636, nc2637, nc2638, 
        nc2639, \B_DOUT_TEMPR6[9] , \B_DOUT_TEMPR6[8] , 
        \B_DOUT_TEMPR6[7] , \B_DOUT_TEMPR6[6] , \B_DOUT_TEMPR6[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[6][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[1] , A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[1] , B_ADDR[13], \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1547 (.A(\B_DOUT_TEMPR56[39] ), .B(\B_DOUT_TEMPR57[39] ), 
        .C(\B_DOUT_TEMPR58[39] ), .D(\B_DOUT_TEMPR59[39] ), .Y(
        OR4_1547_Y));
    OR4 OR4_633 (.A(\A_DOUT_TEMPR16[35] ), .B(\A_DOUT_TEMPR17[35] ), 
        .C(\A_DOUT_TEMPR18[35] ), .D(\A_DOUT_TEMPR19[35] ), .Y(
        OR4_633_Y));
    OR4 OR4_2258 (.A(OR4_778_Y), .B(OR4_2440_Y), .C(OR4_1820_Y), .D(
        OR4_1175_Y), .Y(OR4_2258_Y));
    OR4 OR4_206 (.A(\A_DOUT_TEMPR40[38] ), .B(\A_DOUT_TEMPR41[38] ), 
        .C(\A_DOUT_TEMPR42[38] ), .D(\A_DOUT_TEMPR43[38] ), .Y(
        OR4_206_Y));
    OR4 OR4_25 (.A(\B_DOUT_TEMPR60[39] ), .B(\B_DOUT_TEMPR61[39] ), .C(
        \B_DOUT_TEMPR62[39] ), .D(\B_DOUT_TEMPR63[39] ), .Y(OR4_25_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%101%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R101C4 (
        .A_DOUT({nc2640, nc2641, nc2642, nc2643, nc2644, nc2645, 
        nc2646, nc2647, nc2648, nc2649, nc2650, nc2651, nc2652, nc2653, 
        nc2654, \A_DOUT_TEMPR101[24] , \A_DOUT_TEMPR101[23] , 
        \A_DOUT_TEMPR101[22] , \A_DOUT_TEMPR101[21] , 
        \A_DOUT_TEMPR101[20] }), .B_DOUT({nc2655, nc2656, nc2657, 
        nc2658, nc2659, nc2660, nc2661, nc2662, nc2663, nc2664, nc2665, 
        nc2666, nc2667, nc2668, nc2669, \B_DOUT_TEMPR101[24] , 
        \B_DOUT_TEMPR101[23] , \B_DOUT_TEMPR101[22] , 
        \B_DOUT_TEMPR101[21] , \B_DOUT_TEMPR101[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[101][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR2 OR2_38 (.A(\A_DOUT_TEMPR72[18] ), .B(\A_DOUT_TEMPR73[18] ), .Y(
        OR2_38_Y));
    OR4 OR4_157 (.A(\B_DOUT_TEMPR28[10] ), .B(\B_DOUT_TEMPR29[10] ), 
        .C(\B_DOUT_TEMPR30[10] ), .D(\B_DOUT_TEMPR31[10] ), .Y(
        OR4_157_Y));
    OR4 OR4_1705 (.A(\A_DOUT_TEMPR20[38] ), .B(\A_DOUT_TEMPR21[38] ), 
        .C(\A_DOUT_TEMPR22[38] ), .D(\A_DOUT_TEMPR23[38] ), .Y(
        OR4_1705_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%12%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R12C6 (
        .A_DOUT({nc2670, nc2671, nc2672, nc2673, nc2674, nc2675, 
        nc2676, nc2677, nc2678, nc2679, nc2680, nc2681, nc2682, nc2683, 
        nc2684, \A_DOUT_TEMPR12[34] , \A_DOUT_TEMPR12[33] , 
        \A_DOUT_TEMPR12[32] , \A_DOUT_TEMPR12[31] , 
        \A_DOUT_TEMPR12[30] }), .B_DOUT({nc2685, nc2686, nc2687, 
        nc2688, nc2689, nc2690, nc2691, nc2692, nc2693, nc2694, nc2695, 
        nc2696, nc2697, nc2698, nc2699, \B_DOUT_TEMPR12[34] , 
        \B_DOUT_TEMPR12[33] , \B_DOUT_TEMPR12[32] , 
        \B_DOUT_TEMPR12[31] , \B_DOUT_TEMPR12[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[12][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[32]  (.A(OR4_1050_Y), .B(OR4_1810_Y), .C(OR4_745_Y)
        , .D(OR4_560_Y), .Y(B_DOUT[32]));
    OR4 OR4_979 (.A(\B_DOUT_TEMPR103[20] ), .B(\B_DOUT_TEMPR104[20] ), 
        .C(\B_DOUT_TEMPR105[20] ), .D(\B_DOUT_TEMPR106[20] ), .Y(
        OR4_979_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%19%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R19C0 (
        .A_DOUT({nc2700, nc2701, nc2702, nc2703, nc2704, nc2705, 
        nc2706, nc2707, nc2708, nc2709, nc2710, nc2711, nc2712, nc2713, 
        nc2714, \A_DOUT_TEMPR19[4] , \A_DOUT_TEMPR19[3] , 
        \A_DOUT_TEMPR19[2] , \A_DOUT_TEMPR19[1] , \A_DOUT_TEMPR19[0] })
        , .B_DOUT({nc2715, nc2716, nc2717, nc2718, nc2719, nc2720, 
        nc2721, nc2722, nc2723, nc2724, nc2725, nc2726, nc2727, nc2728, 
        nc2729, \B_DOUT_TEMPR19[4] , \B_DOUT_TEMPR19[3] , 
        \B_DOUT_TEMPR19[2] , \B_DOUT_TEMPR19[1] , \B_DOUT_TEMPR19[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[19][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_799 (.A(\A_DOUT_TEMPR91[32] ), .B(\A_DOUT_TEMPR92[32] ), 
        .C(\A_DOUT_TEMPR93[32] ), .D(\A_DOUT_TEMPR94[32] ), .Y(
        OR4_799_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%117%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R117C4 (
        .A_DOUT({nc2730, nc2731, nc2732, nc2733, nc2734, nc2735, 
        nc2736, nc2737, nc2738, nc2739, nc2740, nc2741, nc2742, nc2743, 
        nc2744, \A_DOUT_TEMPR117[24] , \A_DOUT_TEMPR117[23] , 
        \A_DOUT_TEMPR117[22] , \A_DOUT_TEMPR117[21] , 
        \A_DOUT_TEMPR117[20] }), .B_DOUT({nc2745, nc2746, nc2747, 
        nc2748, nc2749, nc2750, nc2751, nc2752, nc2753, nc2754, nc2755, 
        nc2756, nc2757, nc2758, nc2759, \B_DOUT_TEMPR117[24] , 
        \B_DOUT_TEMPR117[23] , \B_DOUT_TEMPR117[22] , 
        \B_DOUT_TEMPR117[21] , \B_DOUT_TEMPR117[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[117][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_19 (.A(\B_DOUT_TEMPR79[14] ), .B(\B_DOUT_TEMPR80[14] ), .C(
        \B_DOUT_TEMPR81[14] ), .D(\B_DOUT_TEMPR82[14] ), .Y(OR4_19_Y));
    OR4 OR4_563 (.A(\B_DOUT_TEMPR32[13] ), .B(\B_DOUT_TEMPR33[13] ), 
        .C(\B_DOUT_TEMPR34[13] ), .D(\B_DOUT_TEMPR35[13] ), .Y(
        OR4_563_Y));
    OR4 OR4_1563 (.A(\A_DOUT_TEMPR107[34] ), .B(\A_DOUT_TEMPR108[34] ), 
        .C(\A_DOUT_TEMPR109[34] ), .D(\A_DOUT_TEMPR110[34] ), .Y(
        OR4_1563_Y));
    OR4 OR4_2007 (.A(\B_DOUT_TEMPR28[17] ), .B(\B_DOUT_TEMPR29[17] ), 
        .C(\B_DOUT_TEMPR30[17] ), .D(\B_DOUT_TEMPR31[17] ), .Y(
        OR4_2007_Y));
    OR4 OR4_695 (.A(\B_DOUT_TEMPR16[13] ), .B(\B_DOUT_TEMPR17[13] ), 
        .C(\B_DOUT_TEMPR18[13] ), .D(\B_DOUT_TEMPR19[13] ), .Y(
        OR4_695_Y));
    OR4 \OR4_B_DOUT[14]  (.A(OR4_1715_Y), .B(OR4_740_Y), .C(OR4_609_Y), 
        .D(OR4_383_Y), .Y(B_DOUT[14]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%32%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R32C5 (
        .A_DOUT({nc2760, nc2761, nc2762, nc2763, nc2764, nc2765, 
        nc2766, nc2767, nc2768, nc2769, nc2770, nc2771, nc2772, nc2773, 
        nc2774, \A_DOUT_TEMPR32[29] , \A_DOUT_TEMPR32[28] , 
        \A_DOUT_TEMPR32[27] , \A_DOUT_TEMPR32[26] , 
        \A_DOUT_TEMPR32[25] }), .B_DOUT({nc2775, nc2776, nc2777, 
        nc2778, nc2779, nc2780, nc2781, nc2782, nc2783, nc2784, nc2785, 
        nc2786, nc2787, nc2788, nc2789, \B_DOUT_TEMPR32[29] , 
        \B_DOUT_TEMPR32[28] , \B_DOUT_TEMPR32[27] , 
        \B_DOUT_TEMPR32[26] , \B_DOUT_TEMPR32[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[32][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2445 (.A(OR4_1014_Y), .B(OR4_1904_Y), .C(OR4_1547_Y), .D(
        OR4_25_Y), .Y(OR4_2445_Y));
    OR4 OR4_2309 (.A(OR4_888_Y), .B(OR4_1197_Y), .C(OR4_806_Y), .D(
        OR4_1207_Y), .Y(OR4_2309_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%100%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R100C6 (
        .A_DOUT({nc2790, nc2791, nc2792, nc2793, nc2794, nc2795, 
        nc2796, nc2797, nc2798, nc2799, nc2800, nc2801, nc2802, nc2803, 
        nc2804, \A_DOUT_TEMPR100[34] , \A_DOUT_TEMPR100[33] , 
        \A_DOUT_TEMPR100[32] , \A_DOUT_TEMPR100[31] , 
        \A_DOUT_TEMPR100[30] }), .B_DOUT({nc2805, nc2806, nc2807, 
        nc2808, nc2809, nc2810, nc2811, nc2812, nc2813, nc2814, nc2815, 
        nc2816, nc2817, nc2818, nc2819, \B_DOUT_TEMPR100[34] , 
        \B_DOUT_TEMPR100[33] , \B_DOUT_TEMPR100[32] , 
        \B_DOUT_TEMPR100[31] , \B_DOUT_TEMPR100[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[100][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%15%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R15C6 (
        .A_DOUT({nc2820, nc2821, nc2822, nc2823, nc2824, nc2825, 
        nc2826, nc2827, nc2828, nc2829, nc2830, nc2831, nc2832, nc2833, 
        nc2834, \A_DOUT_TEMPR15[34] , \A_DOUT_TEMPR15[33] , 
        \A_DOUT_TEMPR15[32] , \A_DOUT_TEMPR15[31] , 
        \A_DOUT_TEMPR15[30] }), .B_DOUT({nc2835, nc2836, nc2837, 
        nc2838, nc2839, nc2840, nc2841, nc2842, nc2843, nc2844, nc2845, 
        nc2846, nc2847, nc2848, nc2849, \B_DOUT_TEMPR15[34] , 
        \B_DOUT_TEMPR15[33] , \B_DOUT_TEMPR15[32] , 
        \B_DOUT_TEMPR15[31] , \B_DOUT_TEMPR15[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[15][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_483 (.A(\A_DOUT_TEMPR68[18] ), .B(\A_DOUT_TEMPR69[18] ), 
        .C(\A_DOUT_TEMPR70[18] ), .D(\A_DOUT_TEMPR71[18] ), .Y(
        OR4_483_Y));
    OR4 OR4_2977 (.A(\B_DOUT_TEMPR99[24] ), .B(\B_DOUT_TEMPR100[24] ), 
        .C(\B_DOUT_TEMPR101[24] ), .D(\B_DOUT_TEMPR102[24] ), .Y(
        OR4_2977_Y));
    OR4 OR4_2207 (.A(\A_DOUT_TEMPR24[23] ), .B(\A_DOUT_TEMPR25[23] ), 
        .C(\A_DOUT_TEMPR26[23] ), .D(\A_DOUT_TEMPR27[23] ), .Y(
        OR4_2207_Y));
    OR4 OR4_1163 (.A(OR4_311_Y), .B(OR4_1278_Y), .C(OR4_77_Y), .D(
        OR4_2159_Y), .Y(OR4_1163_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%102%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R102C6 (
        .A_DOUT({nc2850, nc2851, nc2852, nc2853, nc2854, nc2855, 
        nc2856, nc2857, nc2858, nc2859, nc2860, nc2861, nc2862, nc2863, 
        nc2864, \A_DOUT_TEMPR102[34] , \A_DOUT_TEMPR102[33] , 
        \A_DOUT_TEMPR102[32] , \A_DOUT_TEMPR102[31] , 
        \A_DOUT_TEMPR102[30] }), .B_DOUT({nc2865, nc2866, nc2867, 
        nc2868, nc2869, nc2870, nc2871, nc2872, nc2873, nc2874, nc2875, 
        nc2876, nc2877, nc2878, nc2879, \B_DOUT_TEMPR102[34] , 
        \B_DOUT_TEMPR102[33] , \B_DOUT_TEMPR102[32] , 
        \B_DOUT_TEMPR102[31] , \B_DOUT_TEMPR102[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[102][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%73%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R73C2 (
        .A_DOUT({nc2880, nc2881, nc2882, nc2883, nc2884, nc2885, 
        nc2886, nc2887, nc2888, nc2889, nc2890, nc2891, nc2892, nc2893, 
        nc2894, \A_DOUT_TEMPR73[14] , \A_DOUT_TEMPR73[13] , 
        \A_DOUT_TEMPR73[12] , \A_DOUT_TEMPR73[11] , 
        \A_DOUT_TEMPR73[10] }), .B_DOUT({nc2895, nc2896, nc2897, 
        nc2898, nc2899, nc2900, nc2901, nc2902, nc2903, nc2904, nc2905, 
        nc2906, nc2907, nc2908, nc2909, \B_DOUT_TEMPR73[14] , 
        \B_DOUT_TEMPR73[13] , \B_DOUT_TEMPR73[12] , 
        \B_DOUT_TEMPR73[11] , \B_DOUT_TEMPR73[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[73][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_299 (.A(\A_DOUT_TEMPR60[2] ), .B(\A_DOUT_TEMPR61[2] ), .C(
        \A_DOUT_TEMPR62[2] ), .D(\A_DOUT_TEMPR63[2] ), .Y(OR4_299_Y));
    OR4 OR4_2290 (.A(\A_DOUT_TEMPR56[2] ), .B(\A_DOUT_TEMPR57[2] ), .C(
        \A_DOUT_TEMPR58[2] ), .D(\A_DOUT_TEMPR59[2] ), .Y(OR4_2290_Y));
    OR4 OR4_1286 (.A(OR4_1148_Y), .B(OR4_2334_Y), .C(OR4_1915_Y), .D(
        OR4_556_Y), .Y(OR4_1286_Y));
    OR4 OR4_2832 (.A(\B_DOUT_TEMPR115[22] ), .B(\B_DOUT_TEMPR116[22] ), 
        .C(\B_DOUT_TEMPR117[22] ), .D(\B_DOUT_TEMPR118[22] ), .Y(
        OR4_2832_Y));
    OR4 OR4_37 (.A(\A_DOUT_TEMPR64[13] ), .B(\A_DOUT_TEMPR65[13] ), .C(
        \A_DOUT_TEMPR66[13] ), .D(\A_DOUT_TEMPR67[13] ), .Y(OR4_37_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%43%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R43C3 (
        .A_DOUT({nc2910, nc2911, nc2912, nc2913, nc2914, nc2915, 
        nc2916, nc2917, nc2918, nc2919, nc2920, nc2921, nc2922, nc2923, 
        nc2924, \A_DOUT_TEMPR43[19] , \A_DOUT_TEMPR43[18] , 
        \A_DOUT_TEMPR43[17] , \A_DOUT_TEMPR43[16] , 
        \A_DOUT_TEMPR43[15] }), .B_DOUT({nc2925, nc2926, nc2927, 
        nc2928, nc2929, nc2930, nc2931, nc2932, nc2933, nc2934, nc2935, 
        nc2936, nc2937, nc2938, nc2939, \B_DOUT_TEMPR43[19] , 
        \B_DOUT_TEMPR43[18] , \B_DOUT_TEMPR43[17] , 
        \B_DOUT_TEMPR43[16] , \B_DOUT_TEMPR43[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[43][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1128 (.A(\A_DOUT_TEMPR91[35] ), .B(\A_DOUT_TEMPR92[35] ), 
        .C(\A_DOUT_TEMPR93[35] ), .D(\A_DOUT_TEMPR94[35] ), .Y(
        OR4_1128_Y));
    OR4 OR4_1062 (.A(\A_DOUT_TEMPR36[17] ), .B(\A_DOUT_TEMPR37[17] ), 
        .C(\A_DOUT_TEMPR38[17] ), .D(\A_DOUT_TEMPR39[17] ), .Y(
        OR4_1062_Y));
    OR4 OR4_3023 (.A(\A_DOUT_TEMPR56[0] ), .B(\A_DOUT_TEMPR57[0] ), .C(
        \A_DOUT_TEMPR58[0] ), .D(\A_DOUT_TEMPR59[0] ), .Y(OR4_3023_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%93%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R93C5 (
        .A_DOUT({nc2940, nc2941, nc2942, nc2943, nc2944, nc2945, 
        nc2946, nc2947, nc2948, nc2949, nc2950, nc2951, nc2952, nc2953, 
        nc2954, \A_DOUT_TEMPR93[29] , \A_DOUT_TEMPR93[28] , 
        \A_DOUT_TEMPR93[27] , \A_DOUT_TEMPR93[26] , 
        \A_DOUT_TEMPR93[25] }), .B_DOUT({nc2955, nc2956, nc2957, 
        nc2958, nc2959, nc2960, nc2961, nc2962, nc2963, nc2964, nc2965, 
        nc2966, nc2967, nc2968, nc2969, \B_DOUT_TEMPR93[29] , 
        \B_DOUT_TEMPR93[28] , \B_DOUT_TEMPR93[27] , 
        \B_DOUT_TEMPR93[26] , \B_DOUT_TEMPR93[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[93][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%32%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R32C1 (
        .A_DOUT({nc2970, nc2971, nc2972, nc2973, nc2974, nc2975, 
        nc2976, nc2977, nc2978, nc2979, nc2980, nc2981, nc2982, nc2983, 
        nc2984, \A_DOUT_TEMPR32[9] , \A_DOUT_TEMPR32[8] , 
        \A_DOUT_TEMPR32[7] , \A_DOUT_TEMPR32[6] , \A_DOUT_TEMPR32[5] })
        , .B_DOUT({nc2985, nc2986, nc2987, nc2988, nc2989, nc2990, 
        nc2991, nc2992, nc2993, nc2994, nc2995, nc2996, nc2997, nc2998, 
        nc2999, \B_DOUT_TEMPR32[9] , \B_DOUT_TEMPR32[8] , 
        \B_DOUT_TEMPR32[7] , \B_DOUT_TEMPR32[6] , \B_DOUT_TEMPR32[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[32][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], 
        A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_793 (.A(\B_DOUT_TEMPR111[33] ), .B(\B_DOUT_TEMPR112[33] ), 
        .C(\B_DOUT_TEMPR113[33] ), .D(\B_DOUT_TEMPR114[33] ), .Y(
        OR4_793_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%65%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R65C2 (
        .A_DOUT({nc3000, nc3001, nc3002, nc3003, nc3004, nc3005, 
        nc3006, nc3007, nc3008, nc3009, nc3010, nc3011, nc3012, nc3013, 
        nc3014, \A_DOUT_TEMPR65[14] , \A_DOUT_TEMPR65[13] , 
        \A_DOUT_TEMPR65[12] , \A_DOUT_TEMPR65[11] , 
        \A_DOUT_TEMPR65[10] }), .B_DOUT({nc3015, nc3016, nc3017, 
        nc3018, nc3019, nc3020, nc3021, nc3022, nc3023, nc3024, nc3025, 
        nc3026, nc3027, nc3028, nc3029, \B_DOUT_TEMPR65[14] , 
        \B_DOUT_TEMPR65[13] , \B_DOUT_TEMPR65[12] , 
        \B_DOUT_TEMPR65[11] , \B_DOUT_TEMPR65[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[65][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2900 (.A(\A_DOUT_TEMPR4[39] ), .B(\A_DOUT_TEMPR5[39] ), .C(
        \A_DOUT_TEMPR6[39] ), .D(\A_DOUT_TEMPR7[39] ), .Y(OR4_2900_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%45%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R45C3 (
        .A_DOUT({nc3030, nc3031, nc3032, nc3033, nc3034, nc3035, 
        nc3036, nc3037, nc3038, nc3039, nc3040, nc3041, nc3042, nc3043, 
        nc3044, \A_DOUT_TEMPR45[19] , \A_DOUT_TEMPR45[18] , 
        \A_DOUT_TEMPR45[17] , \A_DOUT_TEMPR45[16] , 
        \A_DOUT_TEMPR45[15] }), .B_DOUT({nc3045, nc3046, nc3047, 
        nc3048, nc3049, nc3050, nc3051, nc3052, nc3053, nc3054, nc3055, 
        nc3056, nc3057, nc3058, nc3059, \B_DOUT_TEMPR45[19] , 
        \B_DOUT_TEMPR45[18] , \B_DOUT_TEMPR45[17] , 
        \B_DOUT_TEMPR45[16] , \B_DOUT_TEMPR45[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[45][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1832 (.A(\B_DOUT_TEMPR107[25] ), .B(\B_DOUT_TEMPR108[25] ), 
        .C(\B_DOUT_TEMPR109[25] ), .D(\B_DOUT_TEMPR110[25] ), .Y(
        OR4_1832_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_14 (.A(VCC), .B(A_ADDR[18]), .C(
        A_ADDR[17]), .Y(CFG3_14_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%0%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R0C6 (
        .A_DOUT({nc3060, nc3061, nc3062, nc3063, nc3064, nc3065, 
        nc3066, nc3067, nc3068, nc3069, nc3070, nc3071, nc3072, nc3073, 
        nc3074, \A_DOUT_TEMPR0[34] , \A_DOUT_TEMPR0[33] , 
        \A_DOUT_TEMPR0[32] , \A_DOUT_TEMPR0[31] , \A_DOUT_TEMPR0[30] })
        , .B_DOUT({nc3075, nc3076, nc3077, nc3078, nc3079, nc3080, 
        nc3081, nc3082, nc3083, nc3084, nc3085, nc3086, nc3087, nc3088, 
        nc3089, \B_DOUT_TEMPR0[34] , \B_DOUT_TEMPR0[33] , 
        \B_DOUT_TEMPR0[32] , \B_DOUT_TEMPR0[31] , \B_DOUT_TEMPR0[30] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[0][6] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[34], A_DIN[33], A_DIN[32], 
        A_DIN[31], A_DIN[30]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1248 (.A(\B_DOUT_TEMPR64[2] ), .B(\B_DOUT_TEMPR65[2] ), .C(
        \B_DOUT_TEMPR66[2] ), .D(\B_DOUT_TEMPR67[2] ), .Y(OR4_1248_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%26%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R26C3 (
        .A_DOUT({nc3090, nc3091, nc3092, nc3093, nc3094, nc3095, 
        nc3096, nc3097, nc3098, nc3099, nc3100, nc3101, nc3102, nc3103, 
        nc3104, \A_DOUT_TEMPR26[19] , \A_DOUT_TEMPR26[18] , 
        \A_DOUT_TEMPR26[17] , \A_DOUT_TEMPR26[16] , 
        \A_DOUT_TEMPR26[15] }), .B_DOUT({nc3105, nc3106, nc3107, 
        nc3108, nc3109, nc3110, nc3111, nc3112, nc3113, nc3114, nc3115, 
        nc3116, nc3117, nc3118, nc3119, \B_DOUT_TEMPR26[19] , 
        \B_DOUT_TEMPR26[18] , \B_DOUT_TEMPR26[17] , 
        \B_DOUT_TEMPR26[16] , \B_DOUT_TEMPR26[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[26][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[9]  (.A(CFG3_5_Y), .B(CFG3_7_Y), 
        .Y(\BLKX2[9] ));
    OR4 OR4_1957 (.A(\B_DOUT_TEMPR60[36] ), .B(\B_DOUT_TEMPR61[36] ), 
        .C(\B_DOUT_TEMPR62[36] ), .D(\B_DOUT_TEMPR63[36] ), .Y(
        OR4_1957_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%115%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R115C6 (
        .A_DOUT({nc3120, nc3121, nc3122, nc3123, nc3124, nc3125, 
        nc3126, nc3127, nc3128, nc3129, nc3130, nc3131, nc3132, nc3133, 
        nc3134, \A_DOUT_TEMPR115[34] , \A_DOUT_TEMPR115[33] , 
        \A_DOUT_TEMPR115[32] , \A_DOUT_TEMPR115[31] , 
        \A_DOUT_TEMPR115[30] }), .B_DOUT({nc3135, nc3136, nc3137, 
        nc3138, nc3139, nc3140, nc3141, nc3142, nc3143, nc3144, nc3145, 
        nc3146, nc3147, nc3148, nc3149, \B_DOUT_TEMPR115[34] , 
        \B_DOUT_TEMPR115[33] , \B_DOUT_TEMPR115[32] , 
        \B_DOUT_TEMPR115[31] , \B_DOUT_TEMPR115[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[115][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2746 (.A(\B_DOUT_TEMPR91[11] ), .B(\B_DOUT_TEMPR92[11] ), 
        .C(\B_DOUT_TEMPR93[11] ), .D(\B_DOUT_TEMPR94[11] ), .Y(
        OR4_2746_Y));
    OR4 OR4_1823 (.A(\B_DOUT_TEMPR48[10] ), .B(\B_DOUT_TEMPR49[10] ), 
        .C(\B_DOUT_TEMPR50[10] ), .D(\B_DOUT_TEMPR51[10] ), .Y(
        OR4_1823_Y));
    OR4 OR4_614 (.A(OR4_588_Y), .B(OR4_391_Y), .C(OR4_1274_Y), .D(
        OR4_2442_Y), .Y(OR4_614_Y));
    OR4 OR4_298 (.A(\A_DOUT_TEMPR75[11] ), .B(\A_DOUT_TEMPR76[11] ), 
        .C(\A_DOUT_TEMPR77[11] ), .D(\A_DOUT_TEMPR78[11] ), .Y(
        OR4_298_Y));
    OR4 OR4_2870 (.A(OR4_424_Y), .B(OR4_1358_Y), .C(OR4_1019_Y), .D(
        OR4_2483_Y), .Y(OR4_2870_Y));
    OR4 OR4_2396 (.A(\B_DOUT_TEMPR36[16] ), .B(\B_DOUT_TEMPR37[16] ), 
        .C(\B_DOUT_TEMPR38[16] ), .D(\B_DOUT_TEMPR39[16] ), .Y(
        OR4_2396_Y));
    OR4 OR4_2280 (.A(\A_DOUT_TEMPR12[29] ), .B(\A_DOUT_TEMPR13[29] ), 
        .C(\A_DOUT_TEMPR14[29] ), .D(\A_DOUT_TEMPR15[29] ), .Y(
        OR4_2280_Y));
    OR4 OR4_833 (.A(\B_DOUT_TEMPR24[26] ), .B(\B_DOUT_TEMPR25[26] ), 
        .C(\B_DOUT_TEMPR26[26] ), .D(\B_DOUT_TEMPR27[26] ), .Y(
        OR4_833_Y));
    OR4 OR4_909 (.A(OR4_1190_Y), .B(OR4_1004_Y), .C(OR2_28_Y), .D(
        \A_DOUT_TEMPR74[37] ), .Y(OR4_909_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%100%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R100C5 (
        .A_DOUT({nc3150, nc3151, nc3152, nc3153, nc3154, nc3155, 
        nc3156, nc3157, nc3158, nc3159, nc3160, nc3161, nc3162, nc3163, 
        nc3164, \A_DOUT_TEMPR100[29] , \A_DOUT_TEMPR100[28] , 
        \A_DOUT_TEMPR100[27] , \A_DOUT_TEMPR100[26] , 
        \A_DOUT_TEMPR100[25] }), .B_DOUT({nc3165, nc3166, nc3167, 
        nc3168, nc3169, nc3170, nc3171, nc3172, nc3173, nc3174, nc3175, 
        nc3176, nc3177, nc3178, nc3179, \B_DOUT_TEMPR100[29] , 
        \B_DOUT_TEMPR100[28] , \B_DOUT_TEMPR100[27] , 
        \B_DOUT_TEMPR100[26] , \B_DOUT_TEMPR100[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[100][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%79%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R79C4 (
        .A_DOUT({nc3180, nc3181, nc3182, nc3183, nc3184, nc3185, 
        nc3186, nc3187, nc3188, nc3189, nc3190, nc3191, nc3192, nc3193, 
        nc3194, \A_DOUT_TEMPR79[24] , \A_DOUT_TEMPR79[23] , 
        \A_DOUT_TEMPR79[22] , \A_DOUT_TEMPR79[21] , 
        \A_DOUT_TEMPR79[20] }), .B_DOUT({nc3195, nc3196, nc3197, 
        nc3198, nc3199, nc3200, nc3201, nc3202, nc3203, nc3204, nc3205, 
        nc3206, nc3207, nc3208, nc3209, \B_DOUT_TEMPR79[24] , 
        \B_DOUT_TEMPR79[23] , \B_DOUT_TEMPR79[22] , 
        \B_DOUT_TEMPR79[21] , \B_DOUT_TEMPR79[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[79][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2702 (.A(\A_DOUT_TEMPR4[9] ), .B(\A_DOUT_TEMPR5[9] ), .C(
        \A_DOUT_TEMPR6[9] ), .D(\A_DOUT_TEMPR7[9] ), .Y(OR4_2702_Y));
    OR4 OR4_2633 (.A(\A_DOUT_TEMPR107[25] ), .B(\A_DOUT_TEMPR108[25] ), 
        .C(\A_DOUT_TEMPR109[25] ), .D(\A_DOUT_TEMPR110[25] ), .Y(
        OR4_2633_Y));
    OR4 OR4_1729 (.A(\A_DOUT_TEMPR36[39] ), .B(\A_DOUT_TEMPR37[39] ), 
        .C(\A_DOUT_TEMPR38[39] ), .D(\A_DOUT_TEMPR39[39] ), .Y(
        OR4_1729_Y));
    OR4 OR4_2939 (.A(\A_DOUT_TEMPR64[29] ), .B(\A_DOUT_TEMPR65[29] ), 
        .C(\A_DOUT_TEMPR66[29] ), .D(\A_DOUT_TEMPR67[29] ), .Y(
        OR4_2939_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%96%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R96C4 (
        .A_DOUT({nc3210, nc3211, nc3212, nc3213, nc3214, nc3215, 
        nc3216, nc3217, nc3218, nc3219, nc3220, nc3221, nc3222, nc3223, 
        nc3224, \A_DOUT_TEMPR96[24] , \A_DOUT_TEMPR96[23] , 
        \A_DOUT_TEMPR96[22] , \A_DOUT_TEMPR96[21] , 
        \A_DOUT_TEMPR96[20] }), .B_DOUT({nc3225, nc3226, nc3227, 
        nc3228, nc3229, nc3230, nc3231, nc3232, nc3233, nc3234, nc3235, 
        nc3236, nc3237, nc3238, nc3239, \B_DOUT_TEMPR96[24] , 
        \B_DOUT_TEMPR96[23] , \B_DOUT_TEMPR96[22] , 
        \B_DOUT_TEMPR96[21] , \B_DOUT_TEMPR96[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[96][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2874 (.A(\B_DOUT_TEMPR28[5] ), .B(\B_DOUT_TEMPR29[5] ), .C(
        \B_DOUT_TEMPR30[5] ), .D(\B_DOUT_TEMPR31[5] ), .Y(OR4_2874_Y));
    OR4 OR4_428 (.A(\A_DOUT_TEMPR87[22] ), .B(\A_DOUT_TEMPR88[22] ), 
        .C(\A_DOUT_TEMPR89[22] ), .D(\A_DOUT_TEMPR90[22] ), .Y(
        OR4_428_Y));
    OR4 OR4_2226 (.A(\A_DOUT_TEMPR20[3] ), .B(\A_DOUT_TEMPR21[3] ), .C(
        \A_DOUT_TEMPR22[3] ), .D(\A_DOUT_TEMPR23[3] ), .Y(OR4_2226_Y));
    OR4 OR4_1633 (.A(\B_DOUT_TEMPR28[26] ), .B(\B_DOUT_TEMPR29[26] ), 
        .C(\B_DOUT_TEMPR30[26] ), .D(\B_DOUT_TEMPR31[26] ), .Y(
        OR4_1633_Y));
    OR4 OR4_1886 (.A(\B_DOUT_TEMPR52[34] ), .B(\B_DOUT_TEMPR53[34] ), 
        .C(\B_DOUT_TEMPR54[34] ), .D(\B_DOUT_TEMPR55[34] ), .Y(
        OR4_1886_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%4%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R4C1 (
        .A_DOUT({nc3240, nc3241, nc3242, nc3243, nc3244, nc3245, 
        nc3246, nc3247, nc3248, nc3249, nc3250, nc3251, nc3252, nc3253, 
        nc3254, \A_DOUT_TEMPR4[9] , \A_DOUT_TEMPR4[8] , 
        \A_DOUT_TEMPR4[7] , \A_DOUT_TEMPR4[6] , \A_DOUT_TEMPR4[5] }), 
        .B_DOUT({nc3255, nc3256, nc3257, nc3258, nc3259, nc3260, 
        nc3261, nc3262, nc3263, nc3264, nc3265, nc3266, nc3267, nc3268, 
        nc3269, \B_DOUT_TEMPR4[9] , \B_DOUT_TEMPR4[8] , 
        \B_DOUT_TEMPR4[7] , \B_DOUT_TEMPR4[6] , \B_DOUT_TEMPR4[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[4][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[1] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%40%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R40C1 (
        .A_DOUT({nc3270, nc3271, nc3272, nc3273, nc3274, nc3275, 
        nc3276, nc3277, nc3278, nc3279, nc3280, nc3281, nc3282, nc3283, 
        nc3284, \A_DOUT_TEMPR40[9] , \A_DOUT_TEMPR40[8] , 
        \A_DOUT_TEMPR40[7] , \A_DOUT_TEMPR40[6] , \A_DOUT_TEMPR40[5] })
        , .B_DOUT({nc3285, nc3286, nc3287, nc3288, nc3289, nc3290, 
        nc3291, nc3292, nc3293, nc3294, nc3295, nc3296, nc3297, nc3298, 
        nc3299, \B_DOUT_TEMPR40[9] , \B_DOUT_TEMPR40[8] , 
        \B_DOUT_TEMPR40[7] , \B_DOUT_TEMPR40[6] , \B_DOUT_TEMPR40[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[40][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_524 (.A(\B_DOUT_TEMPR32[14] ), .B(\B_DOUT_TEMPR33[14] ), 
        .C(\B_DOUT_TEMPR34[14] ), .D(\B_DOUT_TEMPR35[14] ), .Y(
        OR4_524_Y));
    OR4 OR4_3021 (.A(\A_DOUT_TEMPR8[18] ), .B(\A_DOUT_TEMPR9[18] ), .C(
        \A_DOUT_TEMPR10[18] ), .D(\A_DOUT_TEMPR11[18] ), .Y(OR4_3021_Y)
        );
    OR4 OR4_256 (.A(\A_DOUT_TEMPR24[10] ), .B(\A_DOUT_TEMPR25[10] ), 
        .C(\A_DOUT_TEMPR26[10] ), .D(\A_DOUT_TEMPR27[10] ), .Y(
        OR4_256_Y));
    OR4 OR4_1939 (.A(\A_DOUT_TEMPR0[27] ), .B(\A_DOUT_TEMPR1[27] ), .C(
        \A_DOUT_TEMPR2[27] ), .D(\A_DOUT_TEMPR3[27] ), .Y(OR4_1939_Y));
    OR4 OR4_1850 (.A(\B_DOUT_TEMPR24[36] ), .B(\B_DOUT_TEMPR25[36] ), 
        .C(\B_DOUT_TEMPR26[36] ), .D(\B_DOUT_TEMPR27[36] ), .Y(
        OR4_1850_Y));
    OR4 OR4_1126 (.A(\B_DOUT_TEMPR99[34] ), .B(\B_DOUT_TEMPR100[34] ), 
        .C(\B_DOUT_TEMPR101[34] ), .D(\B_DOUT_TEMPR102[34] ), .Y(
        OR4_1126_Y));
    OR4 OR4_30 (.A(OR4_2113_Y), .B(OR4_368_Y), .C(OR4_83_Y), .D(
        OR4_707_Y), .Y(OR4_30_Y));
    OR4 OR4_2386 (.A(\B_DOUT_TEMPR60[20] ), .B(\B_DOUT_TEMPR61[20] ), 
        .C(\B_DOUT_TEMPR62[20] ), .D(\B_DOUT_TEMPR63[20] ), .Y(
        OR4_2386_Y));
    OR4 OR4_1528 (.A(\A_DOUT_TEMPR68[38] ), .B(\A_DOUT_TEMPR69[38] ), 
        .C(\A_DOUT_TEMPR70[38] ), .D(\A_DOUT_TEMPR71[38] ), .Y(
        OR4_1528_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%95%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R95C5 (
        .A_DOUT({nc3300, nc3301, nc3302, nc3303, nc3304, nc3305, 
        nc3306, nc3307, nc3308, nc3309, nc3310, nc3311, nc3312, nc3313, 
        nc3314, \A_DOUT_TEMPR95[29] , \A_DOUT_TEMPR95[28] , 
        \A_DOUT_TEMPR95[27] , \A_DOUT_TEMPR95[26] , 
        \A_DOUT_TEMPR95[25] }), .B_DOUT({nc3315, nc3316, nc3317, 
        nc3318, nc3319, nc3320, nc3321, nc3322, nc3323, nc3324, nc3325, 
        nc3326, nc3327, nc3328, nc3329, \B_DOUT_TEMPR95[29] , 
        \B_DOUT_TEMPR95[28] , \B_DOUT_TEMPR95[27] , 
        \B_DOUT_TEMPR95[26] , \B_DOUT_TEMPR95[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[95][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_132 (.A(\A_DOUT_TEMPR99[10] ), .B(\A_DOUT_TEMPR100[10] ), 
        .C(\A_DOUT_TEMPR101[10] ), .D(\A_DOUT_TEMPR102[10] ), .Y(
        OR4_132_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%105%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R105C2 (
        .A_DOUT({nc3330, nc3331, nc3332, nc3333, nc3334, nc3335, 
        nc3336, nc3337, nc3338, nc3339, nc3340, nc3341, nc3342, nc3343, 
        nc3344, \A_DOUT_TEMPR105[14] , \A_DOUT_TEMPR105[13] , 
        \A_DOUT_TEMPR105[12] , \A_DOUT_TEMPR105[11] , 
        \A_DOUT_TEMPR105[10] }), .B_DOUT({nc3345, nc3346, nc3347, 
        nc3348, nc3349, nc3350, nc3351, nc3352, nc3353, nc3354, nc3355, 
        nc3356, nc3357, nc3358, nc3359, \B_DOUT_TEMPR105[14] , 
        \B_DOUT_TEMPR105[13] , \B_DOUT_TEMPR105[12] , 
        \B_DOUT_TEMPR105[11] , \B_DOUT_TEMPR105[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[105][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1506 (.A(\B_DOUT_TEMPR64[26] ), .B(\B_DOUT_TEMPR65[26] ), 
        .C(\B_DOUT_TEMPR66[26] ), .D(\B_DOUT_TEMPR67[26] ), .Y(
        OR4_1506_Y));
    OR4 OR4_2602 (.A(\A_DOUT_TEMPR79[25] ), .B(\A_DOUT_TEMPR80[25] ), 
        .C(\A_DOUT_TEMPR81[25] ), .D(\A_DOUT_TEMPR82[25] ), .Y(
        OR4_2602_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%108%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R108C0 (
        .A_DOUT({nc3360, nc3361, nc3362, nc3363, nc3364, nc3365, 
        nc3366, nc3367, nc3368, nc3369, nc3370, nc3371, nc3372, nc3373, 
        nc3374, \A_DOUT_TEMPR108[4] , \A_DOUT_TEMPR108[3] , 
        \A_DOUT_TEMPR108[2] , \A_DOUT_TEMPR108[1] , 
        \A_DOUT_TEMPR108[0] }), .B_DOUT({nc3375, nc3376, nc3377, 
        nc3378, nc3379, nc3380, nc3381, nc3382, nc3383, nc3384, nc3385, 
        nc3386, nc3387, nc3388, nc3389, \B_DOUT_TEMPR108[4] , 
        \B_DOUT_TEMPR108[3] , \B_DOUT_TEMPR108[2] , 
        \B_DOUT_TEMPR108[1] , \B_DOUT_TEMPR108[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[108][0] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[4], 
        B_DIN[3], B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_29 (.A(OR4_1666_Y), .B(OR4_1950_Y), .C(OR4_1515_Y), .D(
        OR4_140_Y), .Y(OR4_29_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%94%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R94C5 (
        .A_DOUT({nc3390, nc3391, nc3392, nc3393, nc3394, nc3395, 
        nc3396, nc3397, nc3398, nc3399, nc3400, nc3401, nc3402, nc3403, 
        nc3404, \A_DOUT_TEMPR94[29] , \A_DOUT_TEMPR94[28] , 
        \A_DOUT_TEMPR94[27] , \A_DOUT_TEMPR94[26] , 
        \A_DOUT_TEMPR94[25] }), .B_DOUT({nc3405, nc3406, nc3407, 
        nc3408, nc3409, nc3410, nc3411, nc3412, nc3413, nc3414, nc3415, 
        nc3416, nc3417, nc3418, nc3419, \B_DOUT_TEMPR94[29] , 
        \B_DOUT_TEMPR94[28] , \B_DOUT_TEMPR94[27] , 
        \B_DOUT_TEMPR94[26] , \B_DOUT_TEMPR94[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[94][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[39]  (.A(OR4_1759_Y), .B(OR4_72_Y), .C(OR4_1748_Y), 
        .D(OR4_579_Y), .Y(B_DOUT[39]));
    OR4 OR4_1854 (.A(\B_DOUT_TEMPR83[10] ), .B(\B_DOUT_TEMPR84[10] ), 
        .C(\B_DOUT_TEMPR85[10] ), .D(\B_DOUT_TEMPR86[10] ), .Y(
        OR4_1854_Y));
    OR4 OR4_1707 (.A(\B_DOUT_TEMPR107[16] ), .B(\B_DOUT_TEMPR108[16] ), 
        .C(\B_DOUT_TEMPR109[16] ), .D(\B_DOUT_TEMPR110[16] ), .Y(
        OR4_1707_Y));
    OR4 OR4_2734 (.A(\A_DOUT_TEMPR79[19] ), .B(\A_DOUT_TEMPR80[19] ), 
        .C(\A_DOUT_TEMPR81[19] ), .D(\A_DOUT_TEMPR82[19] ), .Y(
        OR4_2734_Y));
    OR4 OR4_197 (.A(OR4_794_Y), .B(OR4_1111_Y), .C(OR4_2718_Y), .D(
        OR4_572_Y), .Y(OR4_197_Y));
    OR4 OR4_1270 (.A(\B_DOUT_TEMPR48[31] ), .B(\B_DOUT_TEMPR49[31] ), 
        .C(\B_DOUT_TEMPR50[31] ), .D(\B_DOUT_TEMPR51[31] ), .Y(
        OR4_1270_Y));
    OR4 OR4_1501 (.A(OR4_1495_Y), .B(OR4_2304_Y), .C(OR4_1387_Y), .D(
        OR4_210_Y), .Y(OR4_1501_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%109%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R109C6 (
        .A_DOUT({nc3420, nc3421, nc3422, nc3423, nc3424, nc3425, 
        nc3426, nc3427, nc3428, nc3429, nc3430, nc3431, nc3432, nc3433, 
        nc3434, \A_DOUT_TEMPR109[34] , \A_DOUT_TEMPR109[33] , 
        \A_DOUT_TEMPR109[32] , \A_DOUT_TEMPR109[31] , 
        \A_DOUT_TEMPR109[30] }), .B_DOUT({nc3435, nc3436, nc3437, 
        nc3438, nc3439, nc3440, nc3441, nc3442, nc3443, nc3444, nc3445, 
        nc3446, nc3447, nc3448, nc3449, \B_DOUT_TEMPR109[34] , 
        \B_DOUT_TEMPR109[33] , \B_DOUT_TEMPR109[32] , 
        \B_DOUT_TEMPR109[31] , \B_DOUT_TEMPR109[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[109][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_87 (.A(\A_DOUT_TEMPR115[13] ), .B(\A_DOUT_TEMPR116[13] ), 
        .C(\A_DOUT_TEMPR117[13] ), .D(\A_DOUT_TEMPR118[13] ), .Y(
        OR4_87_Y));
    OR4 OR4_2902 (.A(\A_DOUT_TEMPR44[29] ), .B(\A_DOUT_TEMPR45[29] ), 
        .C(\A_DOUT_TEMPR46[29] ), .D(\A_DOUT_TEMPR47[29] ), .Y(
        OR4_2902_Y));
    OR4 OR4_2431 (.A(OR4_1903_Y), .B(OR4_2974_Y), .C(OR4_1614_Y), .D(
        OR4_22_Y), .Y(OR4_2431_Y));
    OR4 OR4_935 (.A(OR4_2953_Y), .B(OR4_189_Y), .C(OR4_2893_Y), .D(
        OR4_203_Y), .Y(OR4_935_Y));
    OR4 OR4_1734 (.A(OR4_1188_Y), .B(OR4_2676_Y), .C(OR4_195_Y), .D(
        OR4_31_Y), .Y(OR4_1734_Y));
    OR4 OR4_435 (.A(\B_DOUT_TEMPR44[14] ), .B(\B_DOUT_TEMPR45[14] ), 
        .C(\B_DOUT_TEMPR46[14] ), .D(\B_DOUT_TEMPR47[14] ), .Y(
        OR4_435_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%9%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R9C0 (
        .A_DOUT({nc3450, nc3451, nc3452, nc3453, nc3454, nc3455, 
        nc3456, nc3457, nc3458, nc3459, nc3460, nc3461, nc3462, nc3463, 
        nc3464, \A_DOUT_TEMPR9[4] , \A_DOUT_TEMPR9[3] , 
        \A_DOUT_TEMPR9[2] , \A_DOUT_TEMPR9[1] , \A_DOUT_TEMPR9[0] }), 
        .B_DOUT({nc3465, nc3466, nc3467, nc3468, nc3469, nc3470, 
        nc3471, nc3472, nc3473, nc3474, nc3475, nc3476, nc3477, nc3478, 
        nc3479, \B_DOUT_TEMPR9[4] , \B_DOUT_TEMPR9[3] , 
        \B_DOUT_TEMPR9[2] , \B_DOUT_TEMPR9[1] , \B_DOUT_TEMPR9[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[9][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[2] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[2] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1512 (.A(OR4_1740_Y), .B(OR4_332_Y), .C(OR4_2570_Y), .D(
        OR4_1490_Y), .Y(OR4_1512_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[14]  (.A(CFG3_19_Y), .B(
        CFG3_15_Y), .Y(\BLKY2[14] ));
    OR4 OR4_1431 (.A(OR4_2344_Y), .B(OR4_717_Y), .C(OR4_2184_Y), .D(
        OR4_720_Y), .Y(OR4_1431_Y));
    OR4 OR4_2492 (.A(\B_DOUT_TEMPR28[3] ), .B(\B_DOUT_TEMPR29[3] ), .C(
        \B_DOUT_TEMPR30[3] ), .D(\B_DOUT_TEMPR31[3] ), .Y(OR4_2492_Y));
    OR4 OR4_1780 (.A(\B_DOUT_TEMPR16[16] ), .B(\B_DOUT_TEMPR17[16] ), 
        .C(\B_DOUT_TEMPR18[16] ), .D(\B_DOUT_TEMPR19[16] ), .Y(
        OR4_1780_Y));
    OR4 OR4_2826 (.A(\B_DOUT_TEMPR8[26] ), .B(\B_DOUT_TEMPR9[26] ), .C(
        \B_DOUT_TEMPR10[26] ), .D(\B_DOUT_TEMPR11[26] ), .Y(OR4_2826_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%113%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R113C0 (
        .A_DOUT({nc3480, nc3481, nc3482, nc3483, nc3484, nc3485, 
        nc3486, nc3487, nc3488, nc3489, nc3490, nc3491, nc3492, nc3493, 
        nc3494, \A_DOUT_TEMPR113[4] , \A_DOUT_TEMPR113[3] , 
        \A_DOUT_TEMPR113[2] , \A_DOUT_TEMPR113[1] , 
        \A_DOUT_TEMPR113[0] }), .B_DOUT({nc3495, nc3496, nc3497, 
        nc3498, nc3499, nc3500, nc3501, nc3502, nc3503, nc3504, nc3505, 
        nc3506, nc3507, nc3508, nc3509, \B_DOUT_TEMPR113[4] , 
        \B_DOUT_TEMPR113[3] , \B_DOUT_TEMPR113[2] , 
        \B_DOUT_TEMPR113[1] , \B_DOUT_TEMPR113[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[113][0] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[4], 
        B_DIN[3], B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2498 (.A(\B_DOUT_TEMPR107[38] ), .B(\B_DOUT_TEMPR108[38] ), 
        .C(\B_DOUT_TEMPR109[38] ), .D(\B_DOUT_TEMPR110[38] ), .Y(
        OR4_2498_Y));
    OR4 OR4_2112 (.A(\A_DOUT_TEMPR48[27] ), .B(\A_DOUT_TEMPR49[27] ), 
        .C(\A_DOUT_TEMPR50[27] ), .D(\A_DOUT_TEMPR51[27] ), .Y(
        OR4_2112_Y));
    OR4 OR4_1376 (.A(\A_DOUT_TEMPR95[30] ), .B(\A_DOUT_TEMPR96[30] ), 
        .C(\A_DOUT_TEMPR97[30] ), .D(\A_DOUT_TEMPR98[30] ), .Y(
        OR4_1376_Y));
    OR4 OR4_529 (.A(\B_DOUT_TEMPR115[20] ), .B(\B_DOUT_TEMPR116[20] ), 
        .C(\B_DOUT_TEMPR117[20] ), .D(\B_DOUT_TEMPR118[20] ), .Y(
        OR4_529_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%62%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R62C5 (
        .A_DOUT({nc3510, nc3511, nc3512, nc3513, nc3514, nc3515, 
        nc3516, nc3517, nc3518, nc3519, nc3520, nc3521, nc3522, nc3523, 
        nc3524, \A_DOUT_TEMPR62[29] , \A_DOUT_TEMPR62[28] , 
        \A_DOUT_TEMPR62[27] , \A_DOUT_TEMPR62[26] , 
        \A_DOUT_TEMPR62[25] }), .B_DOUT({nc3525, nc3526, nc3527, 
        nc3528, nc3529, nc3530, nc3531, nc3532, nc3533, nc3534, nc3535, 
        nc3536, nc3537, nc3538, nc3539, \B_DOUT_TEMPR62[29] , 
        \B_DOUT_TEMPR62[28] , \B_DOUT_TEMPR62[27] , 
        \B_DOUT_TEMPR62[26] , \B_DOUT_TEMPR62[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[62][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%109%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R109C2 (
        .A_DOUT({nc3540, nc3541, nc3542, nc3543, nc3544, nc3545, 
        nc3546, nc3547, nc3548, nc3549, nc3550, nc3551, nc3552, nc3553, 
        nc3554, \A_DOUT_TEMPR109[14] , \A_DOUT_TEMPR109[13] , 
        \A_DOUT_TEMPR109[12] , \A_DOUT_TEMPR109[11] , 
        \A_DOUT_TEMPR109[10] }), .B_DOUT({nc3555, nc3556, nc3557, 
        nc3558, nc3559, nc3560, nc3561, nc3562, nc3563, nc3564, nc3565, 
        nc3566, nc3567, nc3568, nc3569, \B_DOUT_TEMPR109[14] , 
        \B_DOUT_TEMPR109[13] , \B_DOUT_TEMPR109[12] , 
        \B_DOUT_TEMPR109[11] , \B_DOUT_TEMPR109[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[109][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[29]  (.A(OR4_1163_Y), .B(OR4_831_Y), .C(OR4_690_Y), 
        .D(OR4_2865_Y), .Y(A_DOUT[29]));
    OR4 OR4_448 (.A(\B_DOUT_TEMPR107[14] ), .B(\B_DOUT_TEMPR108[14] ), 
        .C(\B_DOUT_TEMPR109[14] ), .D(\B_DOUT_TEMPR110[14] ), .Y(
        OR4_448_Y));
    OR4 OR4_617 (.A(\B_DOUT_TEMPR28[16] ), .B(\B_DOUT_TEMPR29[16] ), 
        .C(\B_DOUT_TEMPR30[16] ), .D(\B_DOUT_TEMPR31[16] ), .Y(
        OR4_617_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%107%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R107C6 (
        .A_DOUT({nc3570, nc3571, nc3572, nc3573, nc3574, nc3575, 
        nc3576, nc3577, nc3578, nc3579, nc3580, nc3581, nc3582, nc3583, 
        nc3584, \A_DOUT_TEMPR107[34] , \A_DOUT_TEMPR107[33] , 
        \A_DOUT_TEMPR107[32] , \A_DOUT_TEMPR107[31] , 
        \A_DOUT_TEMPR107[30] }), .B_DOUT({nc3585, nc3586, nc3587, 
        nc3588, nc3589, nc3590, nc3591, nc3592, nc3593, nc3594, nc3595, 
        nc3596, nc3597, nc3598, nc3599, \B_DOUT_TEMPR107[34] , 
        \B_DOUT_TEMPR107[33] , \B_DOUT_TEMPR107[32] , 
        \B_DOUT_TEMPR107[31] , \B_DOUT_TEMPR107[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[107][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_544 (.A(\B_DOUT_TEMPR111[24] ), .B(\B_DOUT_TEMPR112[24] ), 
        .C(\B_DOUT_TEMPR113[24] ), .D(\B_DOUT_TEMPR114[24] ), .Y(
        OR4_544_Y));
    OR4 OR4_2547 (.A(OR4_1000_Y), .B(OR4_1928_Y), .C(OR4_1094_Y), .D(
        OR4_1412_Y), .Y(OR4_2547_Y));
    OR4 OR4_2934 (.A(OR4_1125_Y), .B(OR4_126_Y), .C(OR4_329_Y), .D(
        OR4_132_Y), .Y(OR4_2934_Y));
    OR4 OR4_2552 (.A(\B_DOUT_TEMPR24[19] ), .B(\B_DOUT_TEMPR25[19] ), 
        .C(\B_DOUT_TEMPR26[19] ), .D(\B_DOUT_TEMPR27[19] ), .Y(
        OR4_2552_Y));
    OR4 OR4_2482 (.A(OR4_2535_Y), .B(OR4_2337_Y), .C(OR2_53_Y), .D(
        \B_DOUT_TEMPR74[36] ), .Y(OR4_2482_Y));
    OR4 OR4_959 (.A(\A_DOUT_TEMPR40[0] ), .B(\A_DOUT_TEMPR41[0] ), .C(
        \A_DOUT_TEMPR42[0] ), .D(\A_DOUT_TEMPR43[0] ), .Y(OR4_959_Y));
    OR4 OR4_2590 (.A(\B_DOUT_TEMPR91[8] ), .B(\B_DOUT_TEMPR92[8] ), .C(
        \B_DOUT_TEMPR93[8] ), .D(\B_DOUT_TEMPR94[8] ), .Y(OR4_2590_Y));
    OR4 OR4_1934 (.A(OR4_700_Y), .B(OR4_1502_Y), .C(OR2_15_Y), .D(
        \A_DOUT_TEMPR74[28] ), .Y(OR4_1934_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%62%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R62C1 (
        .A_DOUT({nc3600, nc3601, nc3602, nc3603, nc3604, nc3605, 
        nc3606, nc3607, nc3608, nc3609, nc3610, nc3611, nc3612, nc3613, 
        nc3614, \A_DOUT_TEMPR62[9] , \A_DOUT_TEMPR62[8] , 
        \A_DOUT_TEMPR62[7] , \A_DOUT_TEMPR62[6] , \A_DOUT_TEMPR62[5] })
        , .B_DOUT({nc3615, nc3616, nc3617, nc3618, nc3619, nc3620, 
        nc3621, nc3622, nc3623, nc3624, nc3625, nc3626, nc3627, nc3628, 
        nc3629, \B_DOUT_TEMPR62[9] , \B_DOUT_TEMPR62[8] , 
        \B_DOUT_TEMPR62[7] , \B_DOUT_TEMPR62[6] , \B_DOUT_TEMPR62[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[62][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2936 (.A(\A_DOUT_TEMPR32[2] ), .B(\A_DOUT_TEMPR33[2] ), .C(
        \A_DOUT_TEMPR34[2] ), .D(\A_DOUT_TEMPR35[2] ), .Y(OR4_2936_Y));
    OR4 OR4_2488 (.A(\B_DOUT_TEMPR111[29] ), .B(\B_DOUT_TEMPR112[29] ), 
        .C(\B_DOUT_TEMPR113[29] ), .D(\B_DOUT_TEMPR114[29] ), .Y(
        OR4_2488_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%15%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R15C2 (
        .A_DOUT({nc3630, nc3631, nc3632, nc3633, nc3634, nc3635, 
        nc3636, nc3637, nc3638, nc3639, nc3640, nc3641, nc3642, nc3643, 
        nc3644, \A_DOUT_TEMPR15[14] , \A_DOUT_TEMPR15[13] , 
        \A_DOUT_TEMPR15[12] , \A_DOUT_TEMPR15[11] , 
        \A_DOUT_TEMPR15[10] }), .B_DOUT({nc3645, nc3646, nc3647, 
        nc3648, nc3649, nc3650, nc3651, nc3652, nc3653, nc3654, nc3655, 
        nc3656, nc3657, nc3658, nc3659, \B_DOUT_TEMPR15[14] , 
        \B_DOUT_TEMPR15[13] , \B_DOUT_TEMPR15[12] , 
        \B_DOUT_TEMPR15[11] , \B_DOUT_TEMPR15[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[15][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_80 (.A(\B_DOUT_TEMPR79[9] ), .B(\B_DOUT_TEMPR80[9] ), .C(
        \B_DOUT_TEMPR81[9] ), .D(\B_DOUT_TEMPR82[9] ), .Y(OR4_80_Y));
    OR4 OR4_1387 (.A(\A_DOUT_TEMPR111[22] ), .B(\A_DOUT_TEMPR112[22] ), 
        .C(\A_DOUT_TEMPR113[22] ), .D(\A_DOUT_TEMPR114[22] ), .Y(
        OR4_1387_Y));
    OR4 OR4_1282 (.A(\B_DOUT_TEMPR91[31] ), .B(\B_DOUT_TEMPR92[31] ), 
        .C(\B_DOUT_TEMPR93[31] ), .D(\B_DOUT_TEMPR94[31] ), .Y(
        OR4_1282_Y));
    OR4 OR4_1936 (.A(\A_DOUT_TEMPR8[7] ), .B(\A_DOUT_TEMPR9[7] ), .C(
        \A_DOUT_TEMPR10[7] ), .D(\A_DOUT_TEMPR11[7] ), .Y(OR4_1936_Y));
    OR4 OR4_1368 (.A(\A_DOUT_TEMPR87[27] ), .B(\A_DOUT_TEMPR88[27] ), 
        .C(\A_DOUT_TEMPR89[27] ), .D(\A_DOUT_TEMPR90[27] ), .Y(
        OR4_1368_Y));
    OR4 OR4_2720 (.A(\B_DOUT_TEMPR115[4] ), .B(\B_DOUT_TEMPR116[4] ), 
        .C(\B_DOUT_TEMPR117[4] ), .D(\B_DOUT_TEMPR118[4] ), .Y(
        OR4_2720_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%20%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R20C0 (
        .A_DOUT({nc3660, nc3661, nc3662, nc3663, nc3664, nc3665, 
        nc3666, nc3667, nc3668, nc3669, nc3670, nc3671, nc3672, nc3673, 
        nc3674, \A_DOUT_TEMPR20[4] , \A_DOUT_TEMPR20[3] , 
        \A_DOUT_TEMPR20[2] , \A_DOUT_TEMPR20[1] , \A_DOUT_TEMPR20[0] })
        , .B_DOUT({nc3675, nc3676, nc3677, nc3678, nc3679, nc3680, 
        nc3681, nc3682, nc3683, nc3684, nc3685, nc3686, nc3687, nc3688, 
        nc3689, \B_DOUT_TEMPR20[4] , \B_DOUT_TEMPR20[3] , 
        \B_DOUT_TEMPR20[2] , \B_DOUT_TEMPR20[1] , \B_DOUT_TEMPR20[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[20][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%25%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R25C4 (
        .A_DOUT({nc3690, nc3691, nc3692, nc3693, nc3694, nc3695, 
        nc3696, nc3697, nc3698, nc3699, nc3700, nc3701, nc3702, nc3703, 
        nc3704, \A_DOUT_TEMPR25[24] , \A_DOUT_TEMPR25[23] , 
        \A_DOUT_TEMPR25[22] , \A_DOUT_TEMPR25[21] , 
        \A_DOUT_TEMPR25[20] }), .B_DOUT({nc3705, nc3706, nc3707, 
        nc3708, nc3709, nc3710, nc3711, nc3712, nc3713, nc3714, nc3715, 
        nc3716, nc3717, nc3718, nc3719, \B_DOUT_TEMPR25[24] , 
        \B_DOUT_TEMPR25[23] , \B_DOUT_TEMPR25[22] , 
        \B_DOUT_TEMPR25[21] , \B_DOUT_TEMPR25[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[25][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1524 (.A(\B_DOUT_TEMPR79[7] ), .B(\B_DOUT_TEMPR80[7] ), .C(
        \B_DOUT_TEMPR81[7] ), .D(\B_DOUT_TEMPR82[7] ), .Y(OR4_1524_Y));
    OR4 OR4_1010 (.A(OR4_3004_Y), .B(OR4_2825_Y), .C(OR4_2775_Y), .D(
        OR4_336_Y), .Y(OR4_1010_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[16]  (.A(CFG3_11_Y), .B(
        CFG3_21_Y), .Y(\BLKY2[16] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%98%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R98C4 (
        .A_DOUT({nc3720, nc3721, nc3722, nc3723, nc3724, nc3725, 
        nc3726, nc3727, nc3728, nc3729, nc3730, nc3731, nc3732, nc3733, 
        nc3734, \A_DOUT_TEMPR98[24] , \A_DOUT_TEMPR98[23] , 
        \A_DOUT_TEMPR98[22] , \A_DOUT_TEMPR98[21] , 
        \A_DOUT_TEMPR98[20] }), .B_DOUT({nc3735, nc3736, nc3737, 
        nc3738, nc3739, nc3740, nc3741, nc3742, nc3743, nc3744, nc3745, 
        nc3746, nc3747, nc3748, nc3749, \B_DOUT_TEMPR98[24] , 
        \B_DOUT_TEMPR98[23] , \B_DOUT_TEMPR98[22] , 
        \B_DOUT_TEMPR98[21] , \B_DOUT_TEMPR98[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[98][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2409 (.A(\A_DOUT_TEMPR103[20] ), .B(\A_DOUT_TEMPR104[20] ), 
        .C(\A_DOUT_TEMPR105[20] ), .D(\A_DOUT_TEMPR106[20] ), .Y(
        OR4_2409_Y));
    OR4 OR4_2375 (.A(\B_DOUT_TEMPR44[4] ), .B(\B_DOUT_TEMPR45[4] ), .C(
        \B_DOUT_TEMPR46[4] ), .D(\B_DOUT_TEMPR47[4] ), .Y(OR4_2375_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%53%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R53C5 (
        .A_DOUT({nc3750, nc3751, nc3752, nc3753, nc3754, nc3755, 
        nc3756, nc3757, nc3758, nc3759, nc3760, nc3761, nc3762, nc3763, 
        nc3764, \A_DOUT_TEMPR53[29] , \A_DOUT_TEMPR53[28] , 
        \A_DOUT_TEMPR53[27] , \A_DOUT_TEMPR53[26] , 
        \A_DOUT_TEMPR53[25] }), .B_DOUT({nc3765, nc3766, nc3767, 
        nc3768, nc3769, nc3770, nc3771, nc3772, nc3773, nc3774, nc3775, 
        nc3776, nc3777, nc3778, nc3779, \B_DOUT_TEMPR53[29] , 
        \B_DOUT_TEMPR53[28] , \B_DOUT_TEMPR53[27] , 
        \B_DOUT_TEMPR53[26] , \B_DOUT_TEMPR53[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[53][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_35 (.A(OR4_1217_Y), .B(OR4_2226_Y), .C(OR4_939_Y), .D(
        OR4_2324_Y), .Y(OR4_35_Y));
    OR4 OR4_664 (.A(\B_DOUT_TEMPR87[11] ), .B(\B_DOUT_TEMPR88[11] ), 
        .C(\B_DOUT_TEMPR89[11] ), .D(\B_DOUT_TEMPR90[11] ), .Y(
        OR4_664_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%40%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R40C7 (
        .A_DOUT({nc3780, nc3781, nc3782, nc3783, nc3784, nc3785, 
        nc3786, nc3787, nc3788, nc3789, nc3790, nc3791, nc3792, nc3793, 
        nc3794, \A_DOUT_TEMPR40[39] , \A_DOUT_TEMPR40[38] , 
        \A_DOUT_TEMPR40[37] , \A_DOUT_TEMPR40[36] , 
        \A_DOUT_TEMPR40[35] }), .B_DOUT({nc3795, nc3796, nc3797, 
        nc3798, nc3799, nc3800, nc3801, nc3802, nc3803, nc3804, nc3805, 
        nc3806, nc3807, nc3808, nc3809, \B_DOUT_TEMPR40[39] , 
        \B_DOUT_TEMPR40[38] , \B_DOUT_TEMPR40[37] , 
        \B_DOUT_TEMPR40[36] , \B_DOUT_TEMPR40[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[40][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%115%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R115C7 (
        .A_DOUT({nc3810, nc3811, nc3812, nc3813, nc3814, nc3815, 
        nc3816, nc3817, nc3818, nc3819, nc3820, nc3821, nc3822, nc3823, 
        nc3824, \A_DOUT_TEMPR115[39] , \A_DOUT_TEMPR115[38] , 
        \A_DOUT_TEMPR115[37] , \A_DOUT_TEMPR115[36] , 
        \A_DOUT_TEMPR115[35] }), .B_DOUT({nc3825, nc3826, nc3827, 
        nc3828, nc3829, nc3830, nc3831, nc3832, nc3833, nc3834, nc3835, 
        nc3836, nc3837, nc3838, nc3839, \B_DOUT_TEMPR115[39] , 
        \B_DOUT_TEMPR115[38] , \B_DOUT_TEMPR115[37] , 
        \B_DOUT_TEMPR115[36] , \B_DOUT_TEMPR115[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[115][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2580 (.A(\A_DOUT_TEMPR107[33] ), .B(\A_DOUT_TEMPR108[33] ), 
        .C(\A_DOUT_TEMPR109[33] ), .D(\A_DOUT_TEMPR110[33] ), .Y(
        OR4_2580_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%116%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R116C7 (
        .A_DOUT({nc3840, nc3841, nc3842, nc3843, nc3844, nc3845, 
        nc3846, nc3847, nc3848, nc3849, nc3850, nc3851, nc3852, nc3853, 
        nc3854, \A_DOUT_TEMPR116[39] , \A_DOUT_TEMPR116[38] , 
        \A_DOUT_TEMPR116[37] , \A_DOUT_TEMPR116[36] , 
        \A_DOUT_TEMPR116[35] }), .B_DOUT({nc3855, nc3856, nc3857, 
        nc3858, nc3859, nc3860, nc3861, nc3862, nc3863, nc3864, nc3865, 
        nc3866, nc3867, nc3868, nc3869, \B_DOUT_TEMPR116[39] , 
        \B_DOUT_TEMPR116[38] , \B_DOUT_TEMPR116[37] , 
        \B_DOUT_TEMPR116[36] , \B_DOUT_TEMPR116[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[116][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_296 (.A(OR4_321_Y), .B(OR4_1520_Y), .C(OR4_2579_Y), .D(
        OR4_87_Y), .Y(OR4_296_Y));
    OR4 OR4_2260 (.A(\A_DOUT_TEMPR79[22] ), .B(\A_DOUT_TEMPR80[22] ), 
        .C(\A_DOUT_TEMPR81[22] ), .D(\A_DOUT_TEMPR82[22] ), .Y(
        OR4_2260_Y));
    OR4 OR4_217 (.A(\A_DOUT_TEMPR16[38] ), .B(\A_DOUT_TEMPR17[38] ), 
        .C(\A_DOUT_TEMPR18[38] ), .D(\A_DOUT_TEMPR19[38] ), .Y(
        OR4_217_Y));
    OR4 OR4_480 (.A(OR4_403_Y), .B(OR4_211_Y), .C(OR4_150_Y), .D(
        OR4_3039_Y), .Y(OR4_480_Y));
    OR4 OR4_1484 (.A(\A_DOUT_TEMPR20[23] ), .B(\A_DOUT_TEMPR21[23] ), 
        .C(\A_DOUT_TEMPR22[23] ), .D(\A_DOUT_TEMPR23[23] ), .Y(
        OR4_1484_Y));
    OR4 OR4_1472 (.A(\B_DOUT_TEMPR83[38] ), .B(\B_DOUT_TEMPR84[38] ), 
        .C(\B_DOUT_TEMPR85[38] ), .D(\B_DOUT_TEMPR86[38] ), .Y(
        OR4_1472_Y));
    OR4 OR4_1478 (.A(\A_DOUT_TEMPR4[30] ), .B(\A_DOUT_TEMPR5[30] ), .C(
        \A_DOUT_TEMPR6[30] ), .D(\A_DOUT_TEMPR7[30] ), .Y(OR4_1478_Y));
    OR4 OR4_2995 (.A(OR4_1034_Y), .B(OR4_39_Y), .C(OR4_667_Y), .D(
        OR4_2917_Y), .Y(OR4_2995_Y));
    OR4 OR4_1355 (.A(OR4_1959_Y), .B(OR4_3028_Y), .C(OR4_1669_Y), .D(
        OR4_60_Y), .Y(OR4_1355_Y));
    OR4 OR4_1099 (.A(\B_DOUT_TEMPR75[2] ), .B(\B_DOUT_TEMPR76[2] ), .C(
        \B_DOUT_TEMPR77[2] ), .D(\B_DOUT_TEMPR78[2] ), .Y(OR4_1099_Y));
    CFG3 #( .INIT(8'h10) )  CFG3_5 (.A(A_ADDR[16]), .B(A_ADDR[15]), .C(
        A_ADDR[14]), .Y(CFG3_5_Y));
    OR4 OR4_912 (.A(\A_DOUT_TEMPR40[9] ), .B(\A_DOUT_TEMPR41[9] ), .C(
        \A_DOUT_TEMPR42[9] ), .D(\A_DOUT_TEMPR43[9] ), .Y(OR4_912_Y));
    OR4 OR4_549 (.A(\B_DOUT_TEMPR28[23] ), .B(\B_DOUT_TEMPR29[23] ), 
        .C(\B_DOUT_TEMPR30[23] ), .D(\B_DOUT_TEMPR31[23] ), .Y(
        OR4_549_Y));
    OR4 OR4_2327 (.A(\A_DOUT_TEMPR68[14] ), .B(\A_DOUT_TEMPR69[14] ), 
        .C(\A_DOUT_TEMPR70[14] ), .D(\A_DOUT_TEMPR71[14] ), .Y(
        OR4_2327_Y));
    OR4 OR4_2300 (.A(OR4_1993_Y), .B(OR4_2979_Y), .C(OR4_2014_Y), .D(
        OR4_521_Y), .Y(OR4_2300_Y));
    OR4 OR4_1542 (.A(\B_DOUT_TEMPR87[29] ), .B(\B_DOUT_TEMPR88[29] ), 
        .C(\B_DOUT_TEMPR89[29] ), .D(\B_DOUT_TEMPR90[29] ), .Y(
        OR4_1542_Y));
    OR4 OR4_2222 (.A(\A_DOUT_TEMPR68[23] ), .B(\A_DOUT_TEMPR69[23] ), 
        .C(\A_DOUT_TEMPR70[23] ), .D(\A_DOUT_TEMPR71[23] ), .Y(
        OR4_2222_Y));
    OR4 OR4_1221 (.A(\B_DOUT_TEMPR91[4] ), .B(\B_DOUT_TEMPR92[4] ), .C(
        \B_DOUT_TEMPR93[4] ), .D(\B_DOUT_TEMPR94[4] ), .Y(OR4_1221_Y));
    OR4 OR4_2407 (.A(\B_DOUT_TEMPR68[22] ), .B(\B_DOUT_TEMPR69[22] ), 
        .C(\B_DOUT_TEMPR70[22] ), .D(\B_DOUT_TEMPR71[22] ), .Y(
        OR4_2407_Y));
    OR4 OR4_2050 (.A(\A_DOUT_TEMPR103[8] ), .B(\A_DOUT_TEMPR104[8] ), 
        .C(\A_DOUT_TEMPR105[8] ), .D(\A_DOUT_TEMPR106[8] ), .Y(
        OR4_2050_Y));
    OR4 OR4_115 (.A(\A_DOUT_TEMPR87[33] ), .B(\A_DOUT_TEMPR88[33] ), 
        .C(\A_DOUT_TEMPR89[33] ), .D(\A_DOUT_TEMPR90[33] ), .Y(
        OR4_115_Y));
    OR4 OR4_1599 (.A(\A_DOUT_TEMPR20[37] ), .B(\A_DOUT_TEMPR21[37] ), 
        .C(\A_DOUT_TEMPR22[37] ), .D(\A_DOUT_TEMPR23[37] ), .Y(
        OR4_1599_Y));
    OR4 OR4_2248 (.A(OR4_1554_Y), .B(OR4_2545_Y), .C(OR4_174_Y), .D(
        OR4_1848_Y), .Y(OR4_2248_Y));
    OR4 OR4_2699 (.A(OR4_2576_Y), .B(OR4_360_Y), .C(OR4_38_Y), .D(
        OR4_1784_Y), .Y(OR4_2699_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%56%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R56C4 (
        .A_DOUT({nc3870, nc3871, nc3872, nc3873, nc3874, nc3875, 
        nc3876, nc3877, nc3878, nc3879, nc3880, nc3881, nc3882, nc3883, 
        nc3884, \A_DOUT_TEMPR56[24] , \A_DOUT_TEMPR56[23] , 
        \A_DOUT_TEMPR56[22] , \A_DOUT_TEMPR56[21] , 
        \A_DOUT_TEMPR56[20] }), .B_DOUT({nc3885, nc3886, nc3887, 
        nc3888, nc3889, nc3890, nc3891, nc3892, nc3893, nc3894, nc3895, 
        nc3896, nc3897, nc3898, nc3899, \B_DOUT_TEMPR56[24] , 
        \B_DOUT_TEMPR56[23] , \B_DOUT_TEMPR56[22] , 
        \B_DOUT_TEMPR56[21] , \B_DOUT_TEMPR56[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[56][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2366 (.A(\A_DOUT_TEMPR115[23] ), .B(\A_DOUT_TEMPR116[23] ), 
        .C(\A_DOUT_TEMPR117[23] ), .D(\A_DOUT_TEMPR118[23] ), .Y(
        OR4_2366_Y));
    OR4 OR4_910 (.A(\B_DOUT_TEMPR56[0] ), .B(\B_DOUT_TEMPR57[0] ), .C(
        \B_DOUT_TEMPR58[0] ), .D(\B_DOUT_TEMPR59[0] ), .Y(OR4_910_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%109%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R109C4 (
        .A_DOUT({nc3900, nc3901, nc3902, nc3903, nc3904, nc3905, 
        nc3906, nc3907, nc3908, nc3909, nc3910, nc3911, nc3912, nc3913, 
        nc3914, \A_DOUT_TEMPR109[24] , \A_DOUT_TEMPR109[23] , 
        \A_DOUT_TEMPR109[22] , \A_DOUT_TEMPR109[21] , 
        \A_DOUT_TEMPR109[20] }), .B_DOUT({nc3915, nc3916, nc3917, 
        nc3918, nc3919, nc3920, nc3921, nc3922, nc3923, nc3924, nc3925, 
        nc3926, nc3927, nc3928, nc3929, \B_DOUT_TEMPR109[24] , 
        \B_DOUT_TEMPR109[23] , \B_DOUT_TEMPR109[22] , 
        \B_DOUT_TEMPR109[21] , \B_DOUT_TEMPR109[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[109][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%73%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R73C3 (
        .A_DOUT({nc3930, nc3931, nc3932, nc3933, nc3934, nc3935, 
        nc3936, nc3937, nc3938, nc3939, nc3940, nc3941, nc3942, nc3943, 
        nc3944, \A_DOUT_TEMPR73[19] , \A_DOUT_TEMPR73[18] , 
        \A_DOUT_TEMPR73[17] , \A_DOUT_TEMPR73[16] , 
        \A_DOUT_TEMPR73[15] }), .B_DOUT({nc3945, nc3946, nc3947, 
        nc3948, nc3949, nc3950, nc3951, nc3952, nc3953, nc3954, nc3955, 
        nc3956, nc3957, nc3958, nc3959, \B_DOUT_TEMPR73[19] , 
        \B_DOUT_TEMPR73[18] , \B_DOUT_TEMPR73[17] , 
        \B_DOUT_TEMPR73[16] , \B_DOUT_TEMPR73[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[73][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1808 (.A(\B_DOUT_TEMPR75[8] ), .B(\B_DOUT_TEMPR76[8] ), .C(
        \B_DOUT_TEMPR77[8] ), .D(\B_DOUT_TEMPR78[8] ), .Y(OR4_1808_Y));
    OR4 OR4_1465 (.A(\A_DOUT_TEMPR12[23] ), .B(\A_DOUT_TEMPR13[23] ), 
        .C(\A_DOUT_TEMPR14[23] ), .D(\A_DOUT_TEMPR15[23] ), .Y(
        OR4_1465_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%75%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R75C3 (
        .A_DOUT({nc3960, nc3961, nc3962, nc3963, nc3964, nc3965, 
        nc3966, nc3967, nc3968, nc3969, nc3970, nc3971, nc3972, nc3973, 
        nc3974, \A_DOUT_TEMPR75[19] , \A_DOUT_TEMPR75[18] , 
        \A_DOUT_TEMPR75[17] , \A_DOUT_TEMPR75[16] , 
        \A_DOUT_TEMPR75[15] }), .B_DOUT({nc3975, nc3976, nc3977, 
        nc3978, nc3979, nc3980, nc3981, nc3982, nc3983, nc3984, nc3985, 
        nc3986, nc3987, nc3988, nc3989, \B_DOUT_TEMPR75[19] , 
        \B_DOUT_TEMPR75[18] , \B_DOUT_TEMPR75[17] , 
        \B_DOUT_TEMPR75[16] , \B_DOUT_TEMPR75[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[75][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1416 (.A(\B_DOUT_TEMPR8[14] ), .B(\B_DOUT_TEMPR9[14] ), .C(
        \B_DOUT_TEMPR10[14] ), .D(\B_DOUT_TEMPR11[14] ), .Y(OR4_1416_Y)
        );
    OR2 OR2_32 (.A(\B_DOUT_TEMPR72[26] ), .B(\B_DOUT_TEMPR73[26] ), .Y(
        OR2_32_Y));
    OR4 OR4_2219 (.A(OR4_2441_Y), .B(OR4_996_Y), .C(OR4_1797_Y), .D(
        OR4_830_Y), .Y(OR4_2219_Y));
    OR4 OR4_1570 (.A(\B_DOUT_TEMPR52[27] ), .B(\B_DOUT_TEMPR53[27] ), 
        .C(\B_DOUT_TEMPR54[27] ), .D(\B_DOUT_TEMPR55[27] ), .Y(
        OR4_1570_Y));
    OR4 OR4_93 (.A(\A_DOUT_TEMPR56[7] ), .B(\A_DOUT_TEMPR57[7] ), .C(
        \A_DOUT_TEMPR58[7] ), .D(\A_DOUT_TEMPR59[7] ), .Y(OR4_93_Y));
    OR4 OR4_1392 (.A(\A_DOUT_TEMPR83[16] ), .B(\A_DOUT_TEMPR84[16] ), 
        .C(\A_DOUT_TEMPR85[16] ), .D(\A_DOUT_TEMPR86[16] ), .Y(
        OR4_1392_Y));
    OR4 OR4_2985 (.A(\A_DOUT_TEMPR75[1] ), .B(\A_DOUT_TEMPR76[1] ), .C(
        \A_DOUT_TEMPR77[1] ), .D(\A_DOUT_TEMPR78[1] ), .Y(OR4_2985_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%55%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R55C5 (
        .A_DOUT({nc3990, nc3991, nc3992, nc3993, nc3994, nc3995, 
        nc3996, nc3997, nc3998, nc3999, nc4000, nc4001, nc4002, nc4003, 
        nc4004, \A_DOUT_TEMPR55[29] , \A_DOUT_TEMPR55[28] , 
        \A_DOUT_TEMPR55[27] , \A_DOUT_TEMPR55[26] , 
        \A_DOUT_TEMPR55[25] }), .B_DOUT({nc4005, nc4006, nc4007, 
        nc4008, nc4009, nc4010, nc4011, nc4012, nc4013, nc4014, nc4015, 
        nc4016, nc4017, nc4018, nc4019, \B_DOUT_TEMPR55[29] , 
        \B_DOUT_TEMPR55[28] , \B_DOUT_TEMPR55[27] , 
        \B_DOUT_TEMPR55[26] , \B_DOUT_TEMPR55[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[55][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2424 (.A(\A_DOUT_TEMPR99[38] ), .B(\A_DOUT_TEMPR100[38] ), 
        .C(\A_DOUT_TEMPR101[38] ), .D(\A_DOUT_TEMPR102[38] ), .Y(
        OR4_2424_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%54%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R54C5 (
        .A_DOUT({nc4020, nc4021, nc4022, nc4023, nc4024, nc4025, 
        nc4026, nc4027, nc4028, nc4029, nc4030, nc4031, nc4032, nc4033, 
        nc4034, \A_DOUT_TEMPR54[29] , \A_DOUT_TEMPR54[28] , 
        \A_DOUT_TEMPR54[27] , \A_DOUT_TEMPR54[26] , 
        \A_DOUT_TEMPR54[25] }), .B_DOUT({nc4035, nc4036, nc4037, 
        nc4038, nc4039, nc4040, nc4041, nc4042, nc4043, nc4044, nc4045, 
        nc4046, nc4047, nc4048, nc4049, \B_DOUT_TEMPR54[29] , 
        \B_DOUT_TEMPR54[28] , \B_DOUT_TEMPR54[27] , 
        \B_DOUT_TEMPR54[26] , \B_DOUT_TEMPR54[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[54][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_189 (.A(\B_DOUT_TEMPR91[20] ), .B(\B_DOUT_TEMPR92[20] ), 
        .C(\B_DOUT_TEMPR93[20] ), .D(\B_DOUT_TEMPR94[20] ), .Y(
        OR4_189_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%33%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R33C5 (
        .A_DOUT({nc4050, nc4051, nc4052, nc4053, nc4054, nc4055, 
        nc4056, nc4057, nc4058, nc4059, nc4060, nc4061, nc4062, nc4063, 
        nc4064, \A_DOUT_TEMPR33[29] , \A_DOUT_TEMPR33[28] , 
        \A_DOUT_TEMPR33[27] , \A_DOUT_TEMPR33[26] , 
        \A_DOUT_TEMPR33[25] }), .B_DOUT({nc4065, nc4066, nc4067, 
        nc4068, nc4069, nc4070, nc4071, nc4072, nc4073, nc4074, nc4075, 
        nc4076, nc4077, nc4078, nc4079, \B_DOUT_TEMPR33[29] , 
        \B_DOUT_TEMPR33[28] , \B_DOUT_TEMPR33[27] , 
        \B_DOUT_TEMPR33[26] , \B_DOUT_TEMPR33[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[33][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%94%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R94C7 (
        .A_DOUT({nc4080, nc4081, nc4082, nc4083, nc4084, nc4085, 
        nc4086, nc4087, nc4088, nc4089, nc4090, nc4091, nc4092, nc4093, 
        nc4094, \A_DOUT_TEMPR94[39] , \A_DOUT_TEMPR94[38] , 
        \A_DOUT_TEMPR94[37] , \A_DOUT_TEMPR94[36] , 
        \A_DOUT_TEMPR94[35] }), .B_DOUT({nc4095, nc4096, nc4097, 
        nc4098, nc4099, nc4100, nc4101, nc4102, nc4103, nc4104, nc4105, 
        nc4106, nc4107, nc4108, nc4109, \B_DOUT_TEMPR94[39] , 
        \B_DOUT_TEMPR94[38] , \B_DOUT_TEMPR94[37] , 
        \B_DOUT_TEMPR94[36] , \B_DOUT_TEMPR94[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[94][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2689 (.A(OR4_2308_Y), .B(OR4_2950_Y), .C(OR4_1337_Y), .D(
        OR4_2250_Y), .Y(OR4_2689_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%28%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R28C6 (
        .A_DOUT({nc4110, nc4111, nc4112, nc4113, nc4114, nc4115, 
        nc4116, nc4117, nc4118, nc4119, nc4120, nc4121, nc4122, nc4123, 
        nc4124, \A_DOUT_TEMPR28[34] , \A_DOUT_TEMPR28[33] , 
        \A_DOUT_TEMPR28[32] , \A_DOUT_TEMPR28[31] , 
        \A_DOUT_TEMPR28[30] }), .B_DOUT({nc4125, nc4126, nc4127, 
        nc4128, nc4129, nc4130, nc4131, nc4132, nc4133, nc4134, nc4135, 
        nc4136, nc4137, nc4138, nc4139, \B_DOUT_TEMPR28[34] , 
        \B_DOUT_TEMPR28[33] , \B_DOUT_TEMPR28[32] , 
        \B_DOUT_TEMPR28[31] , \B_DOUT_TEMPR28[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[28][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1715 (.A(OR4_238_Y), .B(OR4_1841_Y), .C(OR4_14_Y), .D(
        OR4_2786_Y), .Y(OR4_1715_Y));
    OR4 OR4_85 (.A(\A_DOUT_TEMPR12[14] ), .B(\A_DOUT_TEMPR13[14] ), .C(
        \A_DOUT_TEMPR14[14] ), .D(\A_DOUT_TEMPR15[14] ), .Y(OR4_85_Y));
    OR4 OR4_1766 (.A(\A_DOUT_TEMPR91[9] ), .B(\A_DOUT_TEMPR92[9] ), .C(
        \A_DOUT_TEMPR93[9] ), .D(\A_DOUT_TEMPR94[9] ), .Y(OR4_1766_Y));
    OR4 OR4_1284 (.A(OR4_111_Y), .B(OR4_1120_Y), .C(OR4_1778_Y), .D(
        OR4_413_Y), .Y(OR4_1284_Y));
    OR4 OR4_999 (.A(\A_DOUT_TEMPR91[23] ), .B(\A_DOUT_TEMPR92[23] ), 
        .C(\A_DOUT_TEMPR93[23] ), .D(\A_DOUT_TEMPR94[23] ), .Y(
        OR4_999_Y));
    OR4 OR4_423 (.A(OR4_1699_Y), .B(OR4_229_Y), .C(OR4_1092_Y), .D(
        OR4_85_Y), .Y(OR4_423_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%42%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R42C0 (
        .A_DOUT({nc4140, nc4141, nc4142, nc4143, nc4144, nc4145, 
        nc4146, nc4147, nc4148, nc4149, nc4150, nc4151, nc4152, nc4153, 
        nc4154, \A_DOUT_TEMPR42[4] , \A_DOUT_TEMPR42[3] , 
        \A_DOUT_TEMPR42[2] , \A_DOUT_TEMPR42[1] , \A_DOUT_TEMPR42[0] })
        , .B_DOUT({nc4155, nc4156, nc4157, nc4158, nc4159, nc4160, 
        nc4161, nc4162, nc4163, nc4164, nc4165, nc4166, nc4167, nc4168, 
        nc4169, \B_DOUT_TEMPR42[4] , \B_DOUT_TEMPR42[3] , 
        \B_DOUT_TEMPR42[2] , \B_DOUT_TEMPR42[1] , \B_DOUT_TEMPR42[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[42][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%12%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R12C5 (
        .A_DOUT({nc4170, nc4171, nc4172, nc4173, nc4174, nc4175, 
        nc4176, nc4177, nc4178, nc4179, nc4180, nc4181, nc4182, nc4183, 
        nc4184, \A_DOUT_TEMPR12[29] , \A_DOUT_TEMPR12[28] , 
        \A_DOUT_TEMPR12[27] , \A_DOUT_TEMPR12[26] , 
        \A_DOUT_TEMPR12[25] }), .B_DOUT({nc4185, nc4186, nc4187, 
        nc4188, nc4189, nc4190, nc4191, nc4192, nc4193, nc4194, nc4195, 
        nc4196, nc4197, nc4198, nc4199, \B_DOUT_TEMPR12[29] , 
        \B_DOUT_TEMPR12[28] , \B_DOUT_TEMPR12[27] , 
        \B_DOUT_TEMPR12[26] , \B_DOUT_TEMPR12[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[12][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR2 OR2_27 (.A(\A_DOUT_TEMPR72[22] ), .B(\A_DOUT_TEMPR73[22] ), .Y(
        OR2_27_Y));
    OR4 OR4_2456 (.A(\A_DOUT_TEMPR68[5] ), .B(\A_DOUT_TEMPR69[5] ), .C(
        \A_DOUT_TEMPR70[5] ), .D(\A_DOUT_TEMPR71[5] ), .Y(OR4_2456_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%70%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R70C1 (
        .A_DOUT({nc4200, nc4201, nc4202, nc4203, nc4204, nc4205, 
        nc4206, nc4207, nc4208, nc4209, nc4210, nc4211, nc4212, nc4213, 
        nc4214, \A_DOUT_TEMPR70[9] , \A_DOUT_TEMPR70[8] , 
        \A_DOUT_TEMPR70[7] , \A_DOUT_TEMPR70[6] , \A_DOUT_TEMPR70[5] })
        , .B_DOUT({nc4215, nc4216, nc4217, nc4218, nc4219, nc4220, 
        nc4221, nc4222, nc4223, nc4224, nc4225, nc4226, nc4227, nc4228, 
        nc4229, \B_DOUT_TEMPR70[9] , \B_DOUT_TEMPR70[8] , 
        \B_DOUT_TEMPR70[7] , \B_DOUT_TEMPR70[6] , \B_DOUT_TEMPR70[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[70][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_667 (.A(\A_DOUT_TEMPR40[26] ), .B(\A_DOUT_TEMPR41[26] ), 
        .C(\A_DOUT_TEMPR42[26] ), .D(\A_DOUT_TEMPR43[26] ), .Y(
        OR4_667_Y));
    OR4 OR4_1595 (.A(\A_DOUT_TEMPR95[2] ), .B(\A_DOUT_TEMPR96[2] ), .C(
        \A_DOUT_TEMPR97[2] ), .D(\A_DOUT_TEMPR98[2] ), .Y(OR4_1595_Y));
    OR4 OR4_1040 (.A(\A_DOUT_TEMPR83[9] ), .B(\A_DOUT_TEMPR84[9] ), .C(
        \A_DOUT_TEMPR85[9] ), .D(\A_DOUT_TEMPR86[9] ), .Y(OR4_1040_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%41%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R41C6 (
        .A_DOUT({nc4230, nc4231, nc4232, nc4233, nc4234, nc4235, 
        nc4236, nc4237, nc4238, nc4239, nc4240, nc4241, nc4242, nc4243, 
        nc4244, \A_DOUT_TEMPR41[34] , \A_DOUT_TEMPR41[33] , 
        \A_DOUT_TEMPR41[32] , \A_DOUT_TEMPR41[31] , 
        \A_DOUT_TEMPR41[30] }), .B_DOUT({nc4245, nc4246, nc4247, 
        nc4248, nc4249, nc4250, nc4251, nc4252, nc4253, nc4254, nc4255, 
        nc4256, nc4257, nc4258, nc4259, \B_DOUT_TEMPR41[34] , 
        \B_DOUT_TEMPR41[33] , \B_DOUT_TEMPR41[32] , 
        \B_DOUT_TEMPR41[31] , \B_DOUT_TEMPR41[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[41][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%12%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R12C1 (
        .A_DOUT({nc4260, nc4261, nc4262, nc4263, nc4264, nc4265, 
        nc4266, nc4267, nc4268, nc4269, nc4270, nc4271, nc4272, nc4273, 
        nc4274, \A_DOUT_TEMPR12[9] , \A_DOUT_TEMPR12[8] , 
        \A_DOUT_TEMPR12[7] , \A_DOUT_TEMPR12[6] , \A_DOUT_TEMPR12[5] })
        , .B_DOUT({nc4275, nc4276, nc4277, nc4278, nc4279, nc4280, 
        nc4281, nc4282, nc4283, nc4284, nc4285, nc4286, nc4287, nc4288, 
        nc4289, \B_DOUT_TEMPR12[9] , \B_DOUT_TEMPR12[8] , 
        \B_DOUT_TEMPR12[7] , \B_DOUT_TEMPR12[6] , \B_DOUT_TEMPR12[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[12][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], 
        A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1975 (.A(\A_DOUT_TEMPR79[31] ), .B(\A_DOUT_TEMPR80[31] ), 
        .C(\A_DOUT_TEMPR81[31] ), .D(\A_DOUT_TEMPR82[31] ), .Y(
        OR4_1975_Y));
    OR4 OR4_1708 (.A(\B_DOUT_TEMPR99[10] ), .B(\B_DOUT_TEMPR100[10] ), 
        .C(\B_DOUT_TEMPR101[10] ), .D(\B_DOUT_TEMPR102[10] ), .Y(
        OR4_1708_Y));
    OR4 OR4_1083 (.A(\B_DOUT_TEMPR83[37] ), .B(\B_DOUT_TEMPR84[37] ), 
        .C(\B_DOUT_TEMPR85[37] ), .D(\B_DOUT_TEMPR86[37] ), .Y(
        OR4_1083_Y));
    OR4 OR4_2462 (.A(OR4_2047_Y), .B(OR4_1859_Y), .C(OR2_44_Y), .D(
        \A_DOUT_TEMPR74[32] ), .Y(OR4_2462_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%36%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R36C4 (
        .A_DOUT({nc4290, nc4291, nc4292, nc4293, nc4294, nc4295, 
        nc4296, nc4297, nc4298, nc4299, nc4300, nc4301, nc4302, nc4303, 
        nc4304, \A_DOUT_TEMPR36[24] , \A_DOUT_TEMPR36[23] , 
        \A_DOUT_TEMPR36[22] , \A_DOUT_TEMPR36[21] , 
        \A_DOUT_TEMPR36[20] }), .B_DOUT({nc4305, nc4306, nc4307, 
        nc4308, nc4309, nc4310, nc4311, nc4312, nc4313, nc4314, nc4315, 
        nc4316, nc4317, nc4318, nc4319, \B_DOUT_TEMPR36[24] , 
        \B_DOUT_TEMPR36[23] , \B_DOUT_TEMPR36[22] , 
        \B_DOUT_TEMPR36[21] , \B_DOUT_TEMPR36[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[36][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1681 (.A(\B_DOUT_TEMPR83[32] ), .B(\B_DOUT_TEMPR84[32] ), 
        .C(\B_DOUT_TEMPR85[32] ), .D(\B_DOUT_TEMPR86[32] ), .Y(
        OR4_1681_Y));
    OR4 OR4_39 (.A(\A_DOUT_TEMPR36[26] ), .B(\A_DOUT_TEMPR37[26] ), .C(
        \A_DOUT_TEMPR38[26] ), .D(\A_DOUT_TEMPR39[26] ), .Y(OR4_39_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%3%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R3C3 (
        .A_DOUT({nc4320, nc4321, nc4322, nc4323, nc4324, nc4325, 
        nc4326, nc4327, nc4328, nc4329, nc4330, nc4331, nc4332, nc4333, 
        nc4334, \A_DOUT_TEMPR3[19] , \A_DOUT_TEMPR3[18] , 
        \A_DOUT_TEMPR3[17] , \A_DOUT_TEMPR3[16] , \A_DOUT_TEMPR3[15] })
        , .B_DOUT({nc4335, nc4336, nc4337, nc4338, nc4339, nc4340, 
        nc4341, nc4342, nc4343, nc4344, nc4345, nc4346, nc4347, nc4348, 
        nc4349, \B_DOUT_TEMPR3[19] , \B_DOUT_TEMPR3[18] , 
        \B_DOUT_TEMPR3[17] , \B_DOUT_TEMPR3[16] , \B_DOUT_TEMPR3[15] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[3][3] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[19], A_DIN[18], A_DIN[17], 
        A_DIN[16], A_DIN[15]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2755 (.A(\B_DOUT_TEMPR4[23] ), .B(\B_DOUT_TEMPR5[23] ), .C(
        \B_DOUT_TEMPR6[23] ), .D(\B_DOUT_TEMPR7[23] ), .Y(OR4_2755_Y));
    OR4 OR4_2468 (.A(\B_DOUT_TEMPR8[4] ), .B(\B_DOUT_TEMPR9[4] ), .C(
        \B_DOUT_TEMPR10[4] ), .D(\B_DOUT_TEMPR11[4] ), .Y(OR4_2468_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%116%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R116C0 (
        .A_DOUT({nc4350, nc4351, nc4352, nc4353, nc4354, nc4355, 
        nc4356, nc4357, nc4358, nc4359, nc4360, nc4361, nc4362, nc4363, 
        nc4364, \A_DOUT_TEMPR116[4] , \A_DOUT_TEMPR116[3] , 
        \A_DOUT_TEMPR116[2] , \A_DOUT_TEMPR116[1] , 
        \A_DOUT_TEMPR116[0] }), .B_DOUT({nc4365, nc4366, nc4367, 
        nc4368, nc4369, nc4370, nc4371, nc4372, nc4373, nc4374, nc4375, 
        nc4376, nc4377, nc4378, nc4379, \B_DOUT_TEMPR116[4] , 
        \B_DOUT_TEMPR116[3] , \B_DOUT_TEMPR116[2] , 
        \B_DOUT_TEMPR116[1] , \B_DOUT_TEMPR116[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[116][0] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[4], 
        B_DIN[3], B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_273 (.A(\A_DOUT_TEMPR60[22] ), .B(\A_DOUT_TEMPR61[22] ), 
        .C(\A_DOUT_TEMPR62[22] ), .D(\A_DOUT_TEMPR63[22] ), .Y(
        OR4_273_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%116%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R116C5 (
        .A_DOUT({nc4380, nc4381, nc4382, nc4383, nc4384, nc4385, 
        nc4386, nc4387, nc4388, nc4389, nc4390, nc4391, nc4392, nc4393, 
        nc4394, \A_DOUT_TEMPR116[29] , \A_DOUT_TEMPR116[28] , 
        \A_DOUT_TEMPR116[27] , \A_DOUT_TEMPR116[26] , 
        \A_DOUT_TEMPR116[25] }), .B_DOUT({nc4395, nc4396, nc4397, 
        nc4398, nc4399, nc4400, nc4401, nc4402, nc4403, nc4404, nc4405, 
        nc4406, nc4407, nc4408, nc4409, \B_DOUT_TEMPR116[29] , 
        \B_DOUT_TEMPR116[28] , \B_DOUT_TEMPR116[27] , 
        \B_DOUT_TEMPR116[26] , \B_DOUT_TEMPR116[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[116][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_371 (.A(\A_DOUT_TEMPR87[38] ), .B(\A_DOUT_TEMPR88[38] ), 
        .C(\A_DOUT_TEMPR89[38] ), .D(\A_DOUT_TEMPR90[38] ), .Y(
        OR4_371_Y));
    OR4 OR4_1679 (.A(\A_DOUT_TEMPR52[6] ), .B(\A_DOUT_TEMPR53[6] ), .C(
        \A_DOUT_TEMPR54[6] ), .D(\A_DOUT_TEMPR55[6] ), .Y(OR4_1679_Y));
    OR4 OR4_1783 (.A(\B_DOUT_TEMPR111[10] ), .B(\B_DOUT_TEMPR112[10] ), 
        .C(\B_DOUT_TEMPR113[10] ), .D(\B_DOUT_TEMPR114[10] ), .Y(
        OR4_1783_Y));
    OR4 OR4_875 (.A(\B_DOUT_TEMPR87[2] ), .B(\B_DOUT_TEMPR88[2] ), .C(
        \B_DOUT_TEMPR89[2] ), .D(\B_DOUT_TEMPR90[2] ), .Y(OR4_875_Y));
    OR4 OR4_173 (.A(\B_DOUT_TEMPR36[17] ), .B(\B_DOUT_TEMPR37[17] ), 
        .C(\B_DOUT_TEMPR38[17] ), .D(\B_DOUT_TEMPR39[17] ), .Y(
        OR4_173_Y));
    OR2 OR2_34 (.A(\A_DOUT_TEMPR72[38] ), .B(\A_DOUT_TEMPR73[38] ), .Y(
        OR2_34_Y));
    OR4 OR4_781 (.A(\B_DOUT_TEMPR56[11] ), .B(\B_DOUT_TEMPR57[11] ), 
        .C(\B_DOUT_TEMPR58[11] ), .D(\B_DOUT_TEMPR59[11] ), .Y(
        OR4_781_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%35%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R35C5 (
        .A_DOUT({nc4410, nc4411, nc4412, nc4413, nc4414, nc4415, 
        nc4416, nc4417, nc4418, nc4419, nc4420, nc4421, nc4422, nc4423, 
        nc4424, \A_DOUT_TEMPR35[29] , \A_DOUT_TEMPR35[28] , 
        \A_DOUT_TEMPR35[27] , \A_DOUT_TEMPR35[26] , 
        \A_DOUT_TEMPR35[25] }), .B_DOUT({nc4425, nc4426, nc4427, 
        nc4428, nc4429, nc4430, nc4431, nc4432, nc4433, nc4434, nc4435, 
        nc4436, nc4437, nc4438, nc4439, \B_DOUT_TEMPR35[29] , 
        \B_DOUT_TEMPR35[28] , \B_DOUT_TEMPR35[27] , 
        \B_DOUT_TEMPR35[26] , \B_DOUT_TEMPR35[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[35][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1185 (.A(\B_DOUT_TEMPR0[20] ), .B(\B_DOUT_TEMPR1[20] ), .C(
        \B_DOUT_TEMPR2[20] ), .D(\B_DOUT_TEMPR3[20] ), .Y(OR4_1185_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKX1[0]  (.A(A_ADDR[13]), .Y(
        \BLKX1[0] ));
    OR4 OR4_639 (.A(\A_DOUT_TEMPR75[35] ), .B(\A_DOUT_TEMPR76[35] ), 
        .C(\A_DOUT_TEMPR77[35] ), .D(\A_DOUT_TEMPR78[35] ), .Y(
        OR4_639_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%24%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R24C3 (
        .A_DOUT({nc4440, nc4441, nc4442, nc4443, nc4444, nc4445, 
        nc4446, nc4447, nc4448, nc4449, nc4450, nc4451, nc4452, nc4453, 
        nc4454, \A_DOUT_TEMPR24[19] , \A_DOUT_TEMPR24[18] , 
        \A_DOUT_TEMPR24[17] , \A_DOUT_TEMPR24[16] , 
        \A_DOUT_TEMPR24[15] }), .B_DOUT({nc4455, nc4456, nc4457, 
        nc4458, nc4459, nc4460, nc4461, nc4462, nc4463, nc4464, nc4465, 
        nc4466, nc4467, nc4468, nc4469, \B_DOUT_TEMPR24[19] , 
        \B_DOUT_TEMPR24[18] , \B_DOUT_TEMPR24[17] , 
        \B_DOUT_TEMPR24[16] , \B_DOUT_TEMPR24[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[24][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2224 (.A(OR4_2840_Y), .B(OR4_1288_Y), .C(OR4_1850_Y), .D(
        OR4_1657_Y), .Y(OR4_2224_Y));
    OR4 OR4_2097 (.A(OR4_1073_Y), .B(OR4_2469_Y), .C(OR2_49_Y), .D(
        \A_DOUT_TEMPR74[6] ), .Y(OR4_2097_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%34%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R34C5 (
        .A_DOUT({nc4470, nc4471, nc4472, nc4473, nc4474, nc4475, 
        nc4476, nc4477, nc4478, nc4479, nc4480, nc4481, nc4482, nc4483, 
        nc4484, \A_DOUT_TEMPR34[29] , \A_DOUT_TEMPR34[28] , 
        \A_DOUT_TEMPR34[27] , \A_DOUT_TEMPR34[26] , 
        \A_DOUT_TEMPR34[25] }), .B_DOUT({nc4485, nc4486, nc4487, 
        nc4488, nc4489, nc4490, nc4491, nc4492, nc4493, nc4494, nc4495, 
        nc4496, nc4497, nc4498, nc4499, \B_DOUT_TEMPR34[29] , 
        \B_DOUT_TEMPR34[28] , \B_DOUT_TEMPR34[27] , 
        \B_DOUT_TEMPR34[26] , \B_DOUT_TEMPR34[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[34][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2399 (.A(\A_DOUT_TEMPR12[32] ), .B(\A_DOUT_TEMPR13[32] ), 
        .C(\A_DOUT_TEMPR14[32] ), .D(\A_DOUT_TEMPR15[32] ), .Y(
        OR4_2399_Y));
    OR4 OR4_2297 (.A(\B_DOUT_TEMPR40[28] ), .B(\B_DOUT_TEMPR41[28] ), 
        .C(\B_DOUT_TEMPR42[28] ), .D(\B_DOUT_TEMPR43[28] ), .Y(
        OR4_2297_Y));
    OR4 OR4_267 (.A(\A_DOUT_TEMPR103[0] ), .B(\A_DOUT_TEMPR104[0] ), 
        .C(\A_DOUT_TEMPR105[0] ), .D(\A_DOUT_TEMPR106[0] ), .Y(
        OR4_267_Y));
    OR4 OR4_2560 (.A(OR4_2703_Y), .B(OR4_2498_Y), .C(OR4_2435_Y), .D(
        OR4_1645_Y), .Y(OR4_2560_Y));
    OR4 OR4_1998 (.A(\B_DOUT_TEMPR91[17] ), .B(\B_DOUT_TEMPR92[17] ), 
        .C(\B_DOUT_TEMPR93[17] ), .D(\B_DOUT_TEMPR94[17] ), .Y(
        OR4_1998_Y));
    OR2 OR2_20 (.A(\B_DOUT_TEMPR72[11] ), .B(\B_DOUT_TEMPR73[11] ), .Y(
        OR2_20_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%81%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R81C5 (
        .A_DOUT({nc4500, nc4501, nc4502, nc4503, nc4504, nc4505, 
        nc4506, nc4507, nc4508, nc4509, nc4510, nc4511, nc4512, nc4513, 
        nc4514, \A_DOUT_TEMPR81[29] , \A_DOUT_TEMPR81[28] , 
        \A_DOUT_TEMPR81[27] , \A_DOUT_TEMPR81[26] , 
        \A_DOUT_TEMPR81[25] }), .B_DOUT({nc4515, nc4516, nc4517, 
        nc4518, nc4519, nc4520, nc4521, nc4522, nc4523, nc4524, nc4525, 
        nc4526, nc4527, nc4528, nc4529, \B_DOUT_TEMPR81[29] , 
        \B_DOUT_TEMPR81[28] , \B_DOUT_TEMPR81[27] , 
        \B_DOUT_TEMPR81[26] , \B_DOUT_TEMPR81[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[81][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR2 OR2_68 (.A(\A_DOUT_TEMPR72[10] ), .B(\A_DOUT_TEMPR73[10] ), .Y(
        OR2_68_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%48%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R48C2 (
        .A_DOUT({nc4530, nc4531, nc4532, nc4533, nc4534, nc4535, 
        nc4536, nc4537, nc4538, nc4539, nc4540, nc4541, nc4542, nc4543, 
        nc4544, \A_DOUT_TEMPR48[14] , \A_DOUT_TEMPR48[13] , 
        \A_DOUT_TEMPR48[12] , \A_DOUT_TEMPR48[11] , 
        \A_DOUT_TEMPR48[10] }), .B_DOUT({nc4545, nc4546, nc4547, 
        nc4548, nc4549, nc4550, nc4551, nc4552, nc4553, nc4554, nc4555, 
        nc4556, nc4557, nc4558, nc4559, \B_DOUT_TEMPR48[14] , 
        \B_DOUT_TEMPR48[13] , \B_DOUT_TEMPR48[12] , 
        \B_DOUT_TEMPR48[11] , \B_DOUT_TEMPR48[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[48][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_933 (.A(\A_DOUT_TEMPR20[7] ), .B(\A_DOUT_TEMPR21[7] ), .C(
        \A_DOUT_TEMPR22[7] ), .D(\A_DOUT_TEMPR23[7] ), .Y(OR4_933_Y));
    OR4 OR4_1081 (.A(\B_DOUT_TEMPR56[10] ), .B(\B_DOUT_TEMPR57[10] ), 
        .C(\B_DOUT_TEMPR58[10] ), .D(\B_DOUT_TEMPR59[10] ), .Y(
        OR4_1081_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%58%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R58C4 (
        .A_DOUT({nc4560, nc4561, nc4562, nc4563, nc4564, nc4565, 
        nc4566, nc4567, nc4568, nc4569, nc4570, nc4571, nc4572, nc4573, 
        nc4574, \A_DOUT_TEMPR58[24] , \A_DOUT_TEMPR58[23] , 
        \A_DOUT_TEMPR58[22] , \A_DOUT_TEMPR58[21] , 
        \A_DOUT_TEMPR58[20] }), .B_DOUT({nc4575, nc4576, nc4577, 
        nc4578, nc4579, nc4580, nc4581, nc4582, nc4583, nc4584, nc4585, 
        nc4586, nc4587, nc4588, nc4589, \B_DOUT_TEMPR58[24] , 
        \B_DOUT_TEMPR58[23] , \B_DOUT_TEMPR58[22] , 
        \B_DOUT_TEMPR58[21] , \B_DOUT_TEMPR58[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[58][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2990 (.A(OR4_1838_Y), .B(OR4_2674_Y), .C(OR2_42_Y), .D(
        \A_DOUT_TEMPR74[20] ), .Y(OR4_2990_Y));
    OR4 OR4_1446 (.A(\A_DOUT_TEMPR28[10] ), .B(\A_DOUT_TEMPR29[10] ), 
        .C(\A_DOUT_TEMPR30[10] ), .D(\A_DOUT_TEMPR31[10] ), .Y(
        OR4_1446_Y));
    OR4 OR4_2023 (.A(\B_DOUT_TEMPR24[10] ), .B(\B_DOUT_TEMPR25[10] ), 
        .C(\B_DOUT_TEMPR26[10] ), .D(\B_DOUT_TEMPR27[10] ), .Y(
        OR4_2023_Y));
    OR4 OR4_882 (.A(OR4_223_Y), .B(OR4_1160_Y), .C(OR4_788_Y), .D(
        OR4_2273_Y), .Y(OR4_882_Y));
    OR4 OR4_443 (.A(OR4_2860_Y), .B(OR4_554_Y), .C(OR4_1263_Y), .D(
        OR4_1539_Y), .Y(OR4_443_Y));
    OR2 OR2_18 (.A(\B_DOUT_TEMPR72[31] ), .B(\B_DOUT_TEMPR73[31] ), .Y(
        OR2_18_Y));
    OR4 OR4_772 (.A(\B_DOUT_TEMPR99[13] ), .B(\B_DOUT_TEMPR100[13] ), 
        .C(\B_DOUT_TEMPR101[13] ), .D(\B_DOUT_TEMPR102[13] ), .Y(
        OR4_772_Y));
    OR4 OR4_962 (.A(\B_DOUT_TEMPR68[30] ), .B(\B_DOUT_TEMPR69[30] ), 
        .C(\B_DOUT_TEMPR70[30] ), .D(\B_DOUT_TEMPR71[30] ), .Y(
        OR4_962_Y));
    OR4 OR4_2621 (.A(\A_DOUT_TEMPR24[7] ), .B(\A_DOUT_TEMPR25[7] ), .C(
        \A_DOUT_TEMPR26[7] ), .D(\A_DOUT_TEMPR27[7] ), .Y(OR4_2621_Y));
    OR4 OR4_2087 (.A(OR4_1934_Y), .B(OR4_2126_Y), .C(OR4_2793_Y), .D(
        OR4_1954_Y), .Y(OR4_2087_Y));
    OR4 OR4_165 (.A(\A_DOUT_TEMPR91[7] ), .B(\A_DOUT_TEMPR92[7] ), .C(
        \A_DOUT_TEMPR93[7] ), .D(\A_DOUT_TEMPR94[7] ), .Y(OR4_165_Y));
    OR4 OR4_376 (.A(\A_DOUT_TEMPR28[2] ), .B(\A_DOUT_TEMPR29[2] ), .C(
        \A_DOUT_TEMPR30[2] ), .D(\A_DOUT_TEMPR31[2] ), .Y(OR4_376_Y));
    OR4 OR4_2389 (.A(\A_DOUT_TEMPR75[12] ), .B(\A_DOUT_TEMPR76[12] ), 
        .C(\A_DOUT_TEMPR77[12] ), .D(\A_DOUT_TEMPR78[12] ), .Y(
        OR4_2389_Y));
    OR4 OR4_2723 (.A(\B_DOUT_TEMPR99[16] ), .B(\B_DOUT_TEMPR100[16] ), 
        .C(\B_DOUT_TEMPR101[16] ), .D(\B_DOUT_TEMPR102[16] ), .Y(
        OR4_2723_Y));
    OR4 OR4_203 (.A(\B_DOUT_TEMPR99[20] ), .B(\B_DOUT_TEMPR100[20] ), 
        .C(\B_DOUT_TEMPR101[20] ), .D(\B_DOUT_TEMPR102[20] ), .Y(
        OR4_203_Y));
    OR4 OR4_2287 (.A(\B_DOUT_TEMPR60[33] ), .B(\B_DOUT_TEMPR61[33] ), 
        .C(\B_DOUT_TEMPR62[33] ), .D(\B_DOUT_TEMPR63[33] ), .Y(
        OR4_2287_Y));
    OR4 OR4_2004 (.A(\A_DOUT_TEMPR107[5] ), .B(\A_DOUT_TEMPR108[5] ), 
        .C(\A_DOUT_TEMPR109[5] ), .D(\A_DOUT_TEMPR110[5] ), .Y(
        OR4_2004_Y));
    OR4 OR4_960 (.A(OR4_586_Y), .B(OR4_2135_Y), .C(OR4_2993_Y), .D(
        OR4_2002_Y), .Y(OR4_960_Y));
    OR4 OR4_301 (.A(\A_DOUT_TEMPR83[11] ), .B(\A_DOUT_TEMPR84[11] ), 
        .C(\A_DOUT_TEMPR85[11] ), .D(\A_DOUT_TEMPR86[11] ), .Y(
        OR4_301_Y));
    OR4 OR4_2006 (.A(\A_DOUT_TEMPR16[39] ), .B(\A_DOUT_TEMPR17[39] ), 
        .C(\A_DOUT_TEMPR18[39] ), .D(\A_DOUT_TEMPR19[39] ), .Y(
        OR4_2006_Y));
    OR4 OR4_1516 (.A(\B_DOUT_TEMPR12[37] ), .B(\B_DOUT_TEMPR13[37] ), 
        .C(\B_DOUT_TEMPR14[37] ), .D(\B_DOUT_TEMPR15[37] ), .Y(
        OR4_1516_Y));
    OR4 OR4_2125 (.A(\A_DOUT_TEMPR56[37] ), .B(\A_DOUT_TEMPR57[37] ), 
        .C(\A_DOUT_TEMPR58[37] ), .D(\A_DOUT_TEMPR59[37] ), .Y(
        OR4_2125_Y));
    OR4 OR4_805 (.A(OR4_2933_Y), .B(OR4_1374_Y), .C(OR4_1948_Y), .D(
        OR4_1752_Y), .Y(OR4_805_Y));
    OR4 OR4_1745 (.A(\B_DOUT_TEMPR32[19] ), .B(\B_DOUT_TEMPR33[19] ), 
        .C(\B_DOUT_TEMPR34[19] ), .D(\B_DOUT_TEMPR35[19] ), .Y(
        OR4_1745_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[17]  (.A(CFG3_5_Y), .B(CFG3_3_Y)
        , .Y(\BLKX2[17] ));
    OR4 OR4_103 (.A(\A_DOUT_TEMPR48[31] ), .B(\A_DOUT_TEMPR49[31] ), 
        .C(\A_DOUT_TEMPR50[31] ), .D(\A_DOUT_TEMPR51[31] ), .Y(
        OR4_103_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%48%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R48C3 (
        .A_DOUT({nc4590, nc4591, nc4592, nc4593, nc4594, nc4595, 
        nc4596, nc4597, nc4598, nc4599, nc4600, nc4601, nc4602, nc4603, 
        nc4604, \A_DOUT_TEMPR48[19] , \A_DOUT_TEMPR48[18] , 
        \A_DOUT_TEMPR48[17] , \A_DOUT_TEMPR48[16] , 
        \A_DOUT_TEMPR48[15] }), .B_DOUT({nc4605, nc4606, nc4607, 
        nc4608, nc4609, nc4610, nc4611, nc4612, nc4613, nc4614, nc4615, 
        nc4616, nc4617, nc4618, nc4619, \B_DOUT_TEMPR48[19] , 
        \B_DOUT_TEMPR48[18] , \B_DOUT_TEMPR48[17] , 
        \B_DOUT_TEMPR48[16] , \B_DOUT_TEMPR48[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[48][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1567 (.A(\A_DOUT_TEMPR48[37] ), .B(\A_DOUT_TEMPR49[37] ), 
        .C(\A_DOUT_TEMPR50[37] ), .D(\A_DOUT_TEMPR51[37] ), .Y(
        OR4_1567_Y));
    OR4 OR4_73 (.A(\A_DOUT_TEMPR24[22] ), .B(\A_DOUT_TEMPR25[22] ), .C(
        \A_DOUT_TEMPR26[22] ), .D(\A_DOUT_TEMPR27[22] ), .Y(OR4_73_Y));
    OR4 OR4_577 (.A(\B_DOUT_TEMPR48[5] ), .B(\B_DOUT_TEMPR49[5] ), .C(
        \B_DOUT_TEMPR50[5] ), .D(\B_DOUT_TEMPR51[5] ), .Y(OR4_577_Y));
    OR4 OR4_1717 (.A(OR4_2967_Y), .B(OR4_196_Y), .C(OR4_1803_Y), .D(
        OR4_2750_Y), .Y(OR4_1717_Y));
    OR4 OR4_2792 (.A(\A_DOUT_TEMPR24[16] ), .B(\A_DOUT_TEMPR25[16] ), 
        .C(\A_DOUT_TEMPR26[16] ), .D(\A_DOUT_TEMPR27[16] ), .Y(
        OR4_2792_Y));
    OR4 OR4_2573 (.A(\A_DOUT_TEMPR91[15] ), .B(\A_DOUT_TEMPR92[15] ), 
        .C(\A_DOUT_TEMPR93[15] ), .D(\A_DOUT_TEMPR94[15] ), .Y(
        OR4_2573_Y));
    OR4 OR4_2980 (.A(OR4_2632_Y), .B(OR4_2422_Y), .C(OR4_256_Y), .D(
        OR4_1446_Y), .Y(OR4_2980_Y));
    OR4 OR4_1511 (.A(\B_DOUT_TEMPR20[0] ), .B(\B_DOUT_TEMPR21[0] ), .C(
        \B_DOUT_TEMPR22[0] ), .D(\B_DOUT_TEMPR23[0] ), .Y(OR4_1511_Y));
    OR4 OR4_89 (.A(\A_DOUT_TEMPR8[27] ), .B(\A_DOUT_TEMPR9[27] ), .C(
        \A_DOUT_TEMPR10[27] ), .D(\A_DOUT_TEMPR11[27] ), .Y(OR4_89_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[9]  (.A(CFG3_8_Y), .B(CFG3_15_Y)
        , .Y(\BLKY2[9] ));
    OR4 OR4_1197 (.A(\B_DOUT_TEMPR91[26] ), .B(\B_DOUT_TEMPR92[26] ), 
        .C(\B_DOUT_TEMPR93[26] ), .D(\B_DOUT_TEMPR94[26] ), .Y(
        OR4_1197_Y));
    OR4 OR4_3000 (.A(\A_DOUT_TEMPR12[13] ), .B(\A_DOUT_TEMPR13[13] ), 
        .C(\A_DOUT_TEMPR14[13] ), .D(\A_DOUT_TEMPR15[13] ), .Y(
        OR4_3000_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%44%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R44C1 (
        .A_DOUT({nc4620, nc4621, nc4622, nc4623, nc4624, nc4625, 
        nc4626, nc4627, nc4628, nc4629, nc4630, nc4631, nc4632, nc4633, 
        nc4634, \A_DOUT_TEMPR44[9] , \A_DOUT_TEMPR44[8] , 
        \A_DOUT_TEMPR44[7] , \A_DOUT_TEMPR44[6] , \A_DOUT_TEMPR44[5] })
        , .B_DOUT({nc4635, nc4636, nc4637, nc4638, nc4639, nc4640, 
        nc4641, nc4642, nc4643, nc4644, nc4645, nc4646, nc4647, nc4648, 
        nc4649, \B_DOUT_TEMPR44[9] , \B_DOUT_TEMPR44[8] , 
        \B_DOUT_TEMPR44[7] , \B_DOUT_TEMPR44[6] , \B_DOUT_TEMPR44[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[44][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1694 (.A(\B_DOUT_TEMPR8[23] ), .B(\B_DOUT_TEMPR9[23] ), .C(
        \B_DOUT_TEMPR10[23] ), .D(\B_DOUT_TEMPR11[23] ), .Y(OR4_1694_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%40%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R40C4 (
        .A_DOUT({nc4650, nc4651, nc4652, nc4653, nc4654, nc4655, 
        nc4656, nc4657, nc4658, nc4659, nc4660, nc4661, nc4662, nc4663, 
        nc4664, \A_DOUT_TEMPR40[24] , \A_DOUT_TEMPR40[23] , 
        \A_DOUT_TEMPR40[22] , \A_DOUT_TEMPR40[21] , 
        \A_DOUT_TEMPR40[20] }), .B_DOUT({nc4665, nc4666, nc4667, 
        nc4668, nc4669, nc4670, nc4671, nc4672, nc4673, nc4674, nc4675, 
        nc4676, nc4677, nc4678, nc4679, \B_DOUT_TEMPR40[24] , 
        \B_DOUT_TEMPR40[23] , \B_DOUT_TEMPR40[22] , 
        \B_DOUT_TEMPR40[21] , \B_DOUT_TEMPR40[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[40][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2965 (.A(\B_DOUT_TEMPR95[30] ), .B(\B_DOUT_TEMPR96[30] ), 
        .C(\B_DOUT_TEMPR97[30] ), .D(\B_DOUT_TEMPR98[30] ), .Y(
        OR4_2965_Y));
    OR4 OR4_2173 (.A(OR4_240_Y), .B(OR4_1390_Y), .C(OR4_2877_Y), .D(
        OR4_1392_Y), .Y(OR4_2173_Y));
    OR4 \OR4_B_DOUT[35]  (.A(OR4_156_Y), .B(OR4_394_Y), .C(OR4_1219_Y), 
        .D(OR4_2015_Y), .Y(B_DOUT[35]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%63%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R63C5 (
        .A_DOUT({nc4680, nc4681, nc4682, nc4683, nc4684, nc4685, 
        nc4686, nc4687, nc4688, nc4689, nc4690, nc4691, nc4692, nc4693, 
        nc4694, \A_DOUT_TEMPR63[29] , \A_DOUT_TEMPR63[28] , 
        \A_DOUT_TEMPR63[27] , \A_DOUT_TEMPR63[26] , 
        \A_DOUT_TEMPR63[25] }), .B_DOUT({nc4695, nc4696, nc4697, 
        nc4698, nc4699, nc4700, nc4701, nc4702, nc4703, nc4704, nc4705, 
        nc4706, nc4707, nc4708, nc4709, \B_DOUT_TEMPR63[29] , 
        \B_DOUT_TEMPR63[28] , \B_DOUT_TEMPR63[27] , 
        \B_DOUT_TEMPR63[26] , \B_DOUT_TEMPR63[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[63][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%93%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R93C4 (
        .A_DOUT({nc4710, nc4711, nc4712, nc4713, nc4714, nc4715, 
        nc4716, nc4717, nc4718, nc4719, nc4720, nc4721, nc4722, nc4723, 
        nc4724, \A_DOUT_TEMPR93[24] , \A_DOUT_TEMPR93[23] , 
        \A_DOUT_TEMPR93[22] , \A_DOUT_TEMPR93[21] , 
        \A_DOUT_TEMPR93[20] }), .B_DOUT({nc4725, nc4726, nc4727, 
        nc4728, nc4729, nc4730, nc4731, nc4732, nc4733, nc4734, nc4735, 
        nc4736, nc4737, nc4738, nc4739, \B_DOUT_TEMPR93[24] , 
        \B_DOUT_TEMPR93[23] , \B_DOUT_TEMPR93[22] , 
        \B_DOUT_TEMPR93[21] , \B_DOUT_TEMPR93[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[93][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%70%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R70C7 (
        .A_DOUT({nc4740, nc4741, nc4742, nc4743, nc4744, nc4745, 
        nc4746, nc4747, nc4748, nc4749, nc4750, nc4751, nc4752, nc4753, 
        nc4754, \A_DOUT_TEMPR70[39] , \A_DOUT_TEMPR70[38] , 
        \A_DOUT_TEMPR70[37] , \A_DOUT_TEMPR70[36] , 
        \A_DOUT_TEMPR70[35] }), .B_DOUT({nc4755, nc4756, nc4757, 
        nc4758, nc4759, nc4760, nc4761, nc4762, nc4763, nc4764, nc4765, 
        nc4766, nc4767, nc4768, nc4769, \B_DOUT_TEMPR70[39] , 
        \B_DOUT_TEMPR70[38] , \B_DOUT_TEMPR70[37] , 
        \B_DOUT_TEMPR70[36] , \B_DOUT_TEMPR70[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[70][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2303 (.A(\B_DOUT_TEMPR99[32] ), .B(\B_DOUT_TEMPR100[32] ), 
        .C(\B_DOUT_TEMPR101[32] ), .D(\B_DOUT_TEMPR102[32] ), .Y(
        OR4_2303_Y));
    OR4 OR4_2021 (.A(OR4_342_Y), .B(OR4_1282_Y), .C(OR4_941_Y), .D(
        OR4_2398_Y), .Y(OR4_2021_Y));
    OR4 OR4_2072 (.A(\B_DOUT_TEMPR64[7] ), .B(\B_DOUT_TEMPR65[7] ), .C(
        \B_DOUT_TEMPR66[7] ), .D(\B_DOUT_TEMPR67[7] ), .Y(OR4_2072_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%109%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R109C5 (
        .A_DOUT({nc4770, nc4771, nc4772, nc4773, nc4774, nc4775, 
        nc4776, nc4777, nc4778, nc4779, nc4780, nc4781, nc4782, nc4783, 
        nc4784, \A_DOUT_TEMPR109[29] , \A_DOUT_TEMPR109[28] , 
        \A_DOUT_TEMPR109[27] , \A_DOUT_TEMPR109[26] , 
        \A_DOUT_TEMPR109[25] }), .B_DOUT({nc4785, nc4786, nc4787, 
        nc4788, nc4789, nc4790, nc4791, nc4792, nc4793, nc4794, nc4795, 
        nc4796, nc4797, nc4798, nc4799, \B_DOUT_TEMPR109[29] , 
        \B_DOUT_TEMPR109[28] , \B_DOUT_TEMPR109[27] , 
        \B_DOUT_TEMPR109[26] , \B_DOUT_TEMPR109[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[109][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2669 (.A(OR4_532_Y), .B(OR4_2927_Y), .C(OR4_1770_Y), .D(
        OR4_1749_Y), .Y(OR4_2669_Y));
    OR4 OR4_2542 (.A(\B_DOUT_TEMPR4[34] ), .B(\B_DOUT_TEMPR5[34] ), .C(
        \B_DOUT_TEMPR6[34] ), .D(\B_DOUT_TEMPR7[34] ), .Y(OR4_2542_Y));
    OR4 OR4_1553 (.A(OR4_1995_Y), .B(OR4_1062_Y), .C(OR4_2520_Y), .D(
        OR4_1064_Y), .Y(OR4_1553_Y));
    OR4 OR4_1077 (.A(\B_DOUT_TEMPR68[3] ), .B(\B_DOUT_TEMPR69[3] ), .C(
        \B_DOUT_TEMPR70[3] ), .D(\B_DOUT_TEMPR71[3] ), .Y(OR4_1077_Y));
    OR4 OR4_2692 (.A(OR4_2036_Y), .B(OR4_889_Y), .C(OR4_1568_Y), .D(
        OR4_1864_Y), .Y(OR4_2692_Y));
    OR4 OR4_3039 (.A(\A_DOUT_TEMPR115[37] ), .B(\A_DOUT_TEMPR116[37] ), 
        .C(\A_DOUT_TEMPR117[37] ), .D(\A_DOUT_TEMPR118[37] ), .Y(
        OR4_3039_Y));
    OR4 OR4_2556 (.A(\B_DOUT_TEMPR75[18] ), .B(\B_DOUT_TEMPR76[18] ), 
        .C(\B_DOUT_TEMPR77[18] ), .D(\B_DOUT_TEMPR78[18] ), .Y(
        OR4_2556_Y));
    OR4 OR4_1379 (.A(\A_DOUT_TEMPR95[37] ), .B(\A_DOUT_TEMPR96[37] ), 
        .C(\A_DOUT_TEMPR97[37] ), .D(\A_DOUT_TEMPR98[37] ), .Y(
        OR4_1379_Y));
    OR4 OR4_2782 (.A(\B_DOUT_TEMPR44[13] ), .B(\B_DOUT_TEMPR45[13] ), 
        .C(\B_DOUT_TEMPR46[13] ), .D(\B_DOUT_TEMPR47[13] ), .Y(
        OR4_2782_Y));
    OR4 OR4_702 (.A(\B_DOUT_TEMPR75[32] ), .B(\B_DOUT_TEMPR76[32] ), 
        .C(\B_DOUT_TEMPR77[32] ), .D(\B_DOUT_TEMPR78[32] ), .Y(
        OR4_702_Y));
    OR4 OR4_1277 (.A(\B_DOUT_TEMPR103[8] ), .B(\B_DOUT_TEMPR104[8] ), 
        .C(\B_DOUT_TEMPR105[8] ), .D(\B_DOUT_TEMPR106[8] ), .Y(
        OR4_1277_Y));
    OR4 OR4_2757 (.A(\B_DOUT_TEMPR99[11] ), .B(\B_DOUT_TEMPR100[11] ), 
        .C(\B_DOUT_TEMPR101[11] ), .D(\B_DOUT_TEMPR102[11] ), .Y(
        OR4_2757_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%38%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R38C4 (
        .A_DOUT({nc4800, nc4801, nc4802, nc4803, nc4804, nc4805, 
        nc4806, nc4807, nc4808, nc4809, nc4810, nc4811, nc4812, nc4813, 
        nc4814, \A_DOUT_TEMPR38[24] , \A_DOUT_TEMPR38[23] , 
        \A_DOUT_TEMPR38[22] , \A_DOUT_TEMPR38[21] , 
        \A_DOUT_TEMPR38[20] }), .B_DOUT({nc4815, nc4816, nc4817, 
        nc4818, nc4819, nc4820, nc4821, nc4822, nc4823, nc4824, nc4825, 
        nc4826, nc4827, nc4828, nc4829, \B_DOUT_TEMPR38[24] , 
        \B_DOUT_TEMPR38[23] , \B_DOUT_TEMPR38[22] , 
        \B_DOUT_TEMPR38[21] , \B_DOUT_TEMPR38[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[38][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1153 (.A(\A_DOUT_TEMPR103[9] ), .B(\A_DOUT_TEMPR104[9] ), 
        .C(\A_DOUT_TEMPR105[9] ), .D(\A_DOUT_TEMPR106[9] ), .Y(
        OR4_1153_Y));
    OR4 OR4_306 (.A(OR4_2229_Y), .B(OR4_2717_Y), .C(OR4_282_Y), .D(
        OR4_2516_Y), .Y(OR4_306_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%54%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R54C7 (
        .A_DOUT({nc4830, nc4831, nc4832, nc4833, nc4834, nc4835, 
        nc4836, nc4837, nc4838, nc4839, nc4840, nc4841, nc4842, nc4843, 
        nc4844, \A_DOUT_TEMPR54[39] , \A_DOUT_TEMPR54[38] , 
        \A_DOUT_TEMPR54[37] , \A_DOUT_TEMPR54[36] , 
        \A_DOUT_TEMPR54[35] }), .B_DOUT({nc4845, nc4846, nc4847, 
        nc4848, nc4849, nc4850, nc4851, nc4852, nc4853, nc4854, nc4855, 
        nc4856, nc4857, nc4858, nc4859, \B_DOUT_TEMPR54[39] , 
        \B_DOUT_TEMPR54[38] , \B_DOUT_TEMPR54[37] , 
        \B_DOUT_TEMPR54[36] , \B_DOUT_TEMPR54[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[54][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h20) )  CFG3_15 (.A(B_BLK_EN), .B(B_ADDR[18]), .C(
        B_ADDR[17]), .Y(CFG3_15_Y));
    OR4 OR4_2911 (.A(\A_DOUT_TEMPR75[18] ), .B(\A_DOUT_TEMPR76[18] ), 
        .C(\A_DOUT_TEMPR77[18] ), .D(\A_DOUT_TEMPR78[18] ), .Y(
        OR4_2911_Y));
    OR4 OR4_2551 (.A(\A_DOUT_TEMPR64[24] ), .B(\A_DOUT_TEMPR65[24] ), 
        .C(\A_DOUT_TEMPR66[24] ), .D(\A_DOUT_TEMPR67[24] ), .Y(
        OR4_2551_Y));
    OR4 OR4_2992 (.A(\B_DOUT_TEMPR115[28] ), .B(\B_DOUT_TEMPR116[28] ), 
        .C(\B_DOUT_TEMPR117[28] ), .D(\B_DOUT_TEMPR118[28] ), .Y(
        OR4_2992_Y));
    OR4 OR4_1052 (.A(\B_DOUT_TEMPR107[17] ), .B(\B_DOUT_TEMPR108[17] ), 
        .C(\B_DOUT_TEMPR109[17] ), .D(\B_DOUT_TEMPR110[17] ), .Y(
        OR4_1052_Y));
    OR4 OR4_1970 (.A(\A_DOUT_TEMPR103[19] ), .B(\A_DOUT_TEMPR104[19] ), 
        .C(\A_DOUT_TEMPR105[19] ), .D(\A_DOUT_TEMPR106[19] ), .Y(
        OR4_1970_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%66%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R66C4 (
        .A_DOUT({nc4860, nc4861, nc4862, nc4863, nc4864, nc4865, 
        nc4866, nc4867, nc4868, nc4869, nc4870, nc4871, nc4872, nc4873, 
        nc4874, \A_DOUT_TEMPR66[24] , \A_DOUT_TEMPR66[23] , 
        \A_DOUT_TEMPR66[22] , \A_DOUT_TEMPR66[21] , 
        \A_DOUT_TEMPR66[20] }), .B_DOUT({nc4875, nc4876, nc4877, 
        nc4878, nc4879, nc4880, nc4881, nc4882, nc4883, nc4884, nc4885, 
        nc4886, nc4887, nc4888, nc4889, \B_DOUT_TEMPR66[24] , 
        \B_DOUT_TEMPR66[23] , \B_DOUT_TEMPR66[22] , 
        \B_DOUT_TEMPR66[21] , \B_DOUT_TEMPR66[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[66][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_507 (.A(\A_DOUT_TEMPR87[15] ), .B(\A_DOUT_TEMPR88[15] ), 
        .C(\A_DOUT_TEMPR89[15] ), .D(\A_DOUT_TEMPR90[15] ), .Y(
        OR4_507_Y));
    OR2 OR2_25 (.A(\A_DOUT_TEMPR72[7] ), .B(\A_DOUT_TEMPR73[7] ), .Y(
        OR2_25_Y));
    OR4 OR4_2682 (.A(OR4_2605_Y), .B(OR4_734_Y), .C(OR4_1783_Y), .D(
        OR4_1294_Y), .Y(OR4_2682_Y));
    OR4 OR4_787 (.A(\B_DOUT_TEMPR4[26] ), .B(\B_DOUT_TEMPR5[26] ), .C(
        \B_DOUT_TEMPR6[26] ), .D(\B_DOUT_TEMPR7[26] ), .Y(OR4_787_Y));
    OR4 OR4_1268 (.A(\A_DOUT_TEMPR44[33] ), .B(\A_DOUT_TEMPR45[33] ), 
        .C(\A_DOUT_TEMPR46[33] ), .D(\A_DOUT_TEMPR47[33] ), .Y(
        OR4_1268_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENA[12]  (.A(A_WBYTE_EN[6]), .B(
        A_WEN), .Y(\WBYTEENA[12] ));
    OR4 OR4_1109 (.A(OR4_1264_Y), .B(OR4_262_Y), .C(OR4_476_Y), .D(
        OR4_275_Y), .Y(OR4_1109_Y));
    OR4 OR4_383 (.A(OR4_2288_Y), .B(OR4_448_Y), .C(OR4_1492_Y), .D(
        OR4_582_Y), .Y(OR4_383_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%65%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R65C5 (
        .A_DOUT({nc4890, nc4891, nc4892, nc4893, nc4894, nc4895, 
        nc4896, nc4897, nc4898, nc4899, nc4900, nc4901, nc4902, nc4903, 
        nc4904, \A_DOUT_TEMPR65[29] , \A_DOUT_TEMPR65[28] , 
        \A_DOUT_TEMPR65[27] , \A_DOUT_TEMPR65[26] , 
        \A_DOUT_TEMPR65[25] }), .B_DOUT({nc4905, nc4906, nc4907, 
        nc4908, nc4909, nc4910, nc4911, nc4912, nc4913, nc4914, nc4915, 
        nc4916, nc4917, nc4918, nc4919, \B_DOUT_TEMPR65[29] , 
        \B_DOUT_TEMPR65[28] , \B_DOUT_TEMPR65[27] , 
        \B_DOUT_TEMPR65[26] , \B_DOUT_TEMPR65[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[65][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%91%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R91C4 (
        .A_DOUT({nc4920, nc4921, nc4922, nc4923, nc4924, nc4925, 
        nc4926, nc4927, nc4928, nc4929, nc4930, nc4931, nc4932, nc4933, 
        nc4934, \A_DOUT_TEMPR91[24] , \A_DOUT_TEMPR91[23] , 
        \A_DOUT_TEMPR91[22] , \A_DOUT_TEMPR91[21] , 
        \A_DOUT_TEMPR91[20] }), .B_DOUT({nc4935, nc4936, nc4937, 
        nc4938, nc4939, nc4940, nc4941, nc4942, nc4943, nc4944, nc4945, 
        nc4946, nc4947, nc4948, nc4949, \B_DOUT_TEMPR91[24] , 
        \B_DOUT_TEMPR91[23] , \B_DOUT_TEMPR91[22] , 
        \B_DOUT_TEMPR91[21] , \B_DOUT_TEMPR91[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[91][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[3]  (.A(OR4_2335_Y), .B(OR4_1165_Y), .C(OR4_2771_Y)
        , .D(OR4_2120_Y), .Y(B_DOUT[3]));
    OR4 OR4_2982 (.A(\A_DOUT_TEMPR68[17] ), .B(\A_DOUT_TEMPR69[17] ), 
        .C(\A_DOUT_TEMPR70[17] ), .D(\A_DOUT_TEMPR71[17] ), .Y(
        OR4_2982_Y));
    OR4 OR4_420 (.A(\A_DOUT_TEMPR87[13] ), .B(\A_DOUT_TEMPR88[13] ), 
        .C(\A_DOUT_TEMPR89[13] ), .D(\A_DOUT_TEMPR90[13] ), .Y(
        OR4_420_Y));
    OR4 OR4_788 (.A(\A_DOUT_TEMPR56[30] ), .B(\A_DOUT_TEMPR57[30] ), 
        .C(\A_DOUT_TEMPR58[30] ), .D(\A_DOUT_TEMPR59[30] ), .Y(
        OR4_788_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%64%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R64C5 (
        .A_DOUT({nc4950, nc4951, nc4952, nc4953, nc4954, nc4955, 
        nc4956, nc4957, nc4958, nc4959, nc4960, nc4961, nc4962, nc4963, 
        nc4964, \A_DOUT_TEMPR64[29] , \A_DOUT_TEMPR64[28] , 
        \A_DOUT_TEMPR64[27] , \A_DOUT_TEMPR64[26] , 
        \A_DOUT_TEMPR64[25] }), .B_DOUT({nc4965, nc4966, nc4967, 
        nc4968, nc4969, nc4970, nc4971, nc4972, nc4973, nc4974, nc4975, 
        nc4976, nc4977, nc4978, nc4979, \B_DOUT_TEMPR64[29] , 
        \B_DOUT_TEMPR64[28] , \B_DOUT_TEMPR64[27] , 
        \B_DOUT_TEMPR64[26] , \B_DOUT_TEMPR64[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[64][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1772 (.A(\A_DOUT_TEMPR48[1] ), .B(\A_DOUT_TEMPR49[1] ), .C(
        \A_DOUT_TEMPR50[1] ), .D(\A_DOUT_TEMPR51[1] ), .Y(OR4_1772_Y));
    OR2 OR2_7 (.A(\B_DOUT_TEMPR72[34] ), .B(\B_DOUT_TEMPR73[34] ), .Y(
        OR2_7_Y));
    OR4 OR4_2213 (.A(\B_DOUT_TEMPR83[2] ), .B(\B_DOUT_TEMPR84[2] ), .C(
        \B_DOUT_TEMPR85[2] ), .D(\B_DOUT_TEMPR86[2] ), .Y(OR4_2213_Y));
    OR4 OR4_683 (.A(\A_DOUT_TEMPR75[8] ), .B(\A_DOUT_TEMPR76[8] ), .C(
        \A_DOUT_TEMPR77[8] ), .D(\A_DOUT_TEMPR78[8] ), .Y(OR4_683_Y));
    OR4 OR4_253 (.A(\A_DOUT_TEMPR36[33] ), .B(\A_DOUT_TEMPR37[33] ), 
        .C(\A_DOUT_TEMPR38[33] ), .D(\A_DOUT_TEMPR39[33] ), .Y(
        OR4_253_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%42%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R42C2 (
        .A_DOUT({nc4980, nc4981, nc4982, nc4983, nc4984, nc4985, 
        nc4986, nc4987, nc4988, nc4989, nc4990, nc4991, nc4992, nc4993, 
        nc4994, \A_DOUT_TEMPR42[14] , \A_DOUT_TEMPR42[13] , 
        \A_DOUT_TEMPR42[12] , \A_DOUT_TEMPR42[11] , 
        \A_DOUT_TEMPR42[10] }), .B_DOUT({nc4995, nc4996, nc4997, 
        nc4998, nc4999, nc5000, nc5001, nc5002, nc5003, nc5004, nc5005, 
        nc5006, nc5007, nc5008, nc5009, \B_DOUT_TEMPR42[14] , 
        \B_DOUT_TEMPR42[13] , \B_DOUT_TEMPR42[12] , 
        \B_DOUT_TEMPR42[11] , \B_DOUT_TEMPR42[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[42][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%117%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R117C2 (
        .A_DOUT({nc5010, nc5011, nc5012, nc5013, nc5014, nc5015, 
        nc5016, nc5017, nc5018, nc5019, nc5020, nc5021, nc5022, nc5023, 
        nc5024, \A_DOUT_TEMPR117[14] , \A_DOUT_TEMPR117[13] , 
        \A_DOUT_TEMPR117[12] , \A_DOUT_TEMPR117[11] , 
        \A_DOUT_TEMPR117[10] }), .B_DOUT({nc5025, nc5026, nc5027, 
        nc5028, nc5029, nc5030, nc5031, nc5032, nc5033, nc5034, nc5035, 
        nc5036, nc5037, nc5038, nc5039, \B_DOUT_TEMPR117[14] , 
        \B_DOUT_TEMPR117[13] , \B_DOUT_TEMPR117[12] , 
        \B_DOUT_TEMPR117[11] , \B_DOUT_TEMPR117[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[117][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_351 (.A(\A_DOUT_TEMPR48[5] ), .B(\A_DOUT_TEMPR49[5] ), .C(
        \A_DOUT_TEMPR50[5] ), .D(\A_DOUT_TEMPR51[5] ), .Y(OR4_351_Y));
    OR4 OR4_776 (.A(\A_DOUT_TEMPR79[7] ), .B(\A_DOUT_TEMPR80[7] ), .C(
        \A_DOUT_TEMPR81[7] ), .D(\A_DOUT_TEMPR82[7] ), .Y(OR4_776_Y));
    OR4 OR4_855 (.A(OR4_234_Y), .B(OR4_1178_Y), .C(OR4_803_Y), .D(
        OR4_2287_Y), .Y(OR4_855_Y));
    OR4 OR4_2040 (.A(OR4_1725_Y), .B(OR4_802_Y), .C(OR4_3037_Y), .D(
        OR4_1960_Y), .Y(OR4_2040_Y));
    OR4 OR4_153 (.A(OR4_1573_Y), .B(OR4_1869_Y), .C(OR4_426_Y), .D(
        OR4_1364_Y), .Y(OR4_153_Y));
    OR4 OR4_1546 (.A(OR4_2198_Y), .B(OR4_250_Y), .C(OR4_1844_Y), .D(
        OR4_2248_Y), .Y(OR4_1546_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%22%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R22C6 (
        .A_DOUT({nc5040, nc5041, nc5042, nc5043, nc5044, nc5045, 
        nc5046, nc5047, nc5048, nc5049, nc5050, nc5051, nc5052, nc5053, 
        nc5054, \A_DOUT_TEMPR22[34] , \A_DOUT_TEMPR22[33] , 
        \A_DOUT_TEMPR22[32] , \A_DOUT_TEMPR22[31] , 
        \A_DOUT_TEMPR22[30] }), .B_DOUT({nc5055, nc5056, nc5057, 
        nc5058, nc5059, nc5060, nc5061, nc5062, nc5063, nc5064, nc5065, 
        nc5066, nc5067, nc5068, nc5069, \B_DOUT_TEMPR22[34] , 
        \B_DOUT_TEMPR22[33] , \B_DOUT_TEMPR22[32] , 
        \B_DOUT_TEMPR22[31] , \B_DOUT_TEMPR22[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[22][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%72%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R72C0 (
        .A_DOUT({nc5070, nc5071, nc5072, nc5073, nc5074, nc5075, 
        nc5076, nc5077, nc5078, nc5079, nc5080, nc5081, nc5082, nc5083, 
        nc5084, \A_DOUT_TEMPR72[4] , \A_DOUT_TEMPR72[3] , 
        \A_DOUT_TEMPR72[2] , \A_DOUT_TEMPR72[1] , \A_DOUT_TEMPR72[0] })
        , .B_DOUT({nc5085, nc5086, nc5087, nc5088, nc5089, nc5090, 
        nc5091, nc5092, nc5093, nc5094, nc5095, nc5096, nc5097, nc5098, 
        nc5099, \B_DOUT_TEMPR72[4] , \B_DOUT_TEMPR72[3] , 
        \B_DOUT_TEMPR72[2] , \B_DOUT_TEMPR72[1] , \B_DOUT_TEMPR72[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[72][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%91%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R91C3 (
        .A_DOUT({nc5100, nc5101, nc5102, nc5103, nc5104, nc5105, 
        nc5106, nc5107, nc5108, nc5109, nc5110, nc5111, nc5112, nc5113, 
        nc5114, \A_DOUT_TEMPR91[19] , \A_DOUT_TEMPR91[18] , 
        \A_DOUT_TEMPR91[17] , \A_DOUT_TEMPR91[16] , 
        \A_DOUT_TEMPR91[15] }), .B_DOUT({nc5115, nc5116, nc5117, 
        nc5118, nc5119, nc5120, nc5121, nc5122, nc5123, nc5124, nc5125, 
        nc5126, nc5127, nc5128, nc5129, \B_DOUT_TEMPR91[19] , 
        \B_DOUT_TEMPR91[18] , \B_DOUT_TEMPR91[17] , 
        \B_DOUT_TEMPR91[16] , \B_DOUT_TEMPR91[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[91][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1747 (.A(\A_DOUT_TEMPR79[10] ), .B(\A_DOUT_TEMPR80[10] ), 
        .C(\A_DOUT_TEMPR81[10] ), .D(\A_DOUT_TEMPR82[10] ), .Y(
        OR4_1747_Y));
    OR4 OR4_436 (.A(\B_DOUT_TEMPR0[39] ), .B(\B_DOUT_TEMPR1[39] ), .C(
        \B_DOUT_TEMPR2[39] ), .D(\B_DOUT_TEMPR3[39] ), .Y(OR4_436_Y));
    OR4 OR4_1541 (.A(OR4_1215_Y), .B(OR4_1794_Y), .C(OR4_184_Y), .D(
        OR4_1161_Y), .Y(OR4_1541_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%34%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R34C7 (
        .A_DOUT({nc5130, nc5131, nc5132, nc5133, nc5134, nc5135, 
        nc5136, nc5137, nc5138, nc5139, nc5140, nc5141, nc5142, nc5143, 
        nc5144, \A_DOUT_TEMPR34[39] , \A_DOUT_TEMPR34[38] , 
        \A_DOUT_TEMPR34[37] , \A_DOUT_TEMPR34[36] , 
        \A_DOUT_TEMPR34[35] }), .B_DOUT({nc5145, nc5146, nc5147, 
        nc5148, nc5149, nc5150, nc5151, nc5152, nc5153, nc5154, nc5155, 
        nc5156, nc5157, nc5158, nc5159, \B_DOUT_TEMPR34[39] , 
        \B_DOUT_TEMPR34[38] , \B_DOUT_TEMPR34[37] , 
        \B_DOUT_TEMPR34[36] , \B_DOUT_TEMPR34[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[34][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%29%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R29C0 (
        .A_DOUT({nc5160, nc5161, nc5162, nc5163, nc5164, nc5165, 
        nc5166, nc5167, nc5168, nc5169, nc5170, nc5171, nc5172, nc5173, 
        nc5174, \A_DOUT_TEMPR29[4] , \A_DOUT_TEMPR29[3] , 
        \A_DOUT_TEMPR29[2] , \A_DOUT_TEMPR29[1] , \A_DOUT_TEMPR29[0] })
        , .B_DOUT({nc5175, nc5176, nc5177, nc5178, nc5179, nc5180, 
        nc5181, nc5182, nc5183, nc5184, nc5185, nc5186, nc5187, nc5188, 
        nc5189, \B_DOUT_TEMPR29[4] , \B_DOUT_TEMPR29[3] , 
        \B_DOUT_TEMPR29[2] , \B_DOUT_TEMPR29[1] , \B_DOUT_TEMPR29[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[29][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1672 (.A(\A_DOUT_TEMPR24[25] ), .B(\A_DOUT_TEMPR25[25] ), 
        .C(\A_DOUT_TEMPR26[25] ), .D(\A_DOUT_TEMPR27[25] ), .Y(
        OR4_1672_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%86%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R86C3 (
        .A_DOUT({nc5190, nc5191, nc5192, nc5193, nc5194, nc5195, 
        nc5196, nc5197, nc5198, nc5199, nc5200, nc5201, nc5202, nc5203, 
        nc5204, \A_DOUT_TEMPR86[19] , \A_DOUT_TEMPR86[18] , 
        \A_DOUT_TEMPR86[17] , \A_DOUT_TEMPR86[16] , 
        \A_DOUT_TEMPR86[15] }), .B_DOUT({nc5205, nc5206, nc5207, 
        nc5208, nc5209, nc5210, nc5211, nc5212, nc5213, nc5214, nc5215, 
        nc5216, nc5217, nc5218, nc5219, \B_DOUT_TEMPR86[19] , 
        \B_DOUT_TEMPR86[18] , \B_DOUT_TEMPR86[17] , 
        \B_DOUT_TEMPR86[16] , \B_DOUT_TEMPR86[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[86][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%71%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R71C6 (
        .A_DOUT({nc5220, nc5221, nc5222, nc5223, nc5224, nc5225, 
        nc5226, nc5227, nc5228, nc5229, nc5230, nc5231, nc5232, nc5233, 
        nc5234, \A_DOUT_TEMPR71[34] , \A_DOUT_TEMPR71[33] , 
        \A_DOUT_TEMPR71[32] , \A_DOUT_TEMPR71[31] , 
        \A_DOUT_TEMPR71[30] }), .B_DOUT({nc5235, nc5236, nc5237, 
        nc5238, nc5239, nc5240, nc5241, nc5242, nc5243, nc5244, nc5245, 
        nc5246, nc5247, nc5248, nc5249, \B_DOUT_TEMPR71[34] , 
        \B_DOUT_TEMPR71[33] , \B_DOUT_TEMPR71[32] , 
        \B_DOUT_TEMPR71[31] , \B_DOUT_TEMPR71[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[71][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1690 (.A(OR4_202_Y), .B(OR4_1221_Y), .C(OR4_1887_Y), .D(
        OR4_513_Y), .Y(OR4_1690_Y));
    OR4 OR4_2067 (.A(\B_DOUT_TEMPR28[25] ), .B(\B_DOUT_TEMPR29[25] ), 
        .C(\B_DOUT_TEMPR30[25] ), .D(\B_DOUT_TEMPR31[25] ), .Y(
        OR4_2067_Y));
    OR4 OR4_2499 (.A(\A_DOUT_TEMPR32[10] ), .B(\A_DOUT_TEMPR33[10] ), 
        .C(\A_DOUT_TEMPR34[10] ), .D(\A_DOUT_TEMPR35[10] ), .Y(
        OR4_2499_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%43%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R43C1 (
        .A_DOUT({nc5250, nc5251, nc5252, nc5253, nc5254, nc5255, 
        nc5256, nc5257, nc5258, nc5259, nc5260, nc5261, nc5262, nc5263, 
        nc5264, \A_DOUT_TEMPR43[9] , \A_DOUT_TEMPR43[8] , 
        \A_DOUT_TEMPR43[7] , \A_DOUT_TEMPR43[6] , \A_DOUT_TEMPR43[5] })
        , .B_DOUT({nc5265, nc5266, nc5267, nc5268, nc5269, nc5270, 
        nc5271, nc5272, nc5273, nc5274, nc5275, nc5276, nc5277, nc5278, 
        nc5279, \B_DOUT_TEMPR43[9] , \B_DOUT_TEMPR43[8] , 
        \B_DOUT_TEMPR43[7] , \B_DOUT_TEMPR43[6] , \B_DOUT_TEMPR43[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[43][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2369 (.A(\B_DOUT_TEMPR99[36] ), .B(\B_DOUT_TEMPR100[36] ), 
        .C(\B_DOUT_TEMPR101[36] ), .D(\B_DOUT_TEMPR102[36] ), .Y(
        OR4_2369_Y));
    OR4 OR4_1972 (.A(\A_DOUT_TEMPR28[27] ), .B(\A_DOUT_TEMPR29[27] ), 
        .C(\A_DOUT_TEMPR30[27] ), .D(\A_DOUT_TEMPR31[27] ), .Y(
        OR4_1972_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%25%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R25C6 (
        .A_DOUT({nc5280, nc5281, nc5282, nc5283, nc5284, nc5285, 
        nc5286, nc5287, nc5288, nc5289, nc5290, nc5291, nc5292, nc5293, 
        nc5294, \A_DOUT_TEMPR25[34] , \A_DOUT_TEMPR25[33] , 
        \A_DOUT_TEMPR25[32] , \A_DOUT_TEMPR25[31] , 
        \A_DOUT_TEMPR25[30] }), .B_DOUT({nc5295, nc5296, nc5297, 
        nc5298, nc5299, nc5300, nc5301, nc5302, nc5303, nc5304, nc5305, 
        nc5306, nc5307, nc5308, nc5309, \B_DOUT_TEMPR25[34] , 
        \B_DOUT_TEMPR25[33] , \B_DOUT_TEMPR25[32] , 
        \B_DOUT_TEMPR25[31] , \B_DOUT_TEMPR25[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[25][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2267 (.A(\A_DOUT_TEMPR111[32] ), .B(\A_DOUT_TEMPR112[32] ), 
        .C(\A_DOUT_TEMPR113[32] ), .D(\A_DOUT_TEMPR114[32] ), .Y(
        OR4_2267_Y));
    OR4 OR4_1098 (.A(OR4_2216_Y), .B(OR4_1247_Y), .C(OR4_2734_Y), .D(
        OR4_1250_Y), .Y(OR4_1098_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%110%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R110C1 (
        .A_DOUT({nc5310, nc5311, nc5312, nc5313, nc5314, nc5315, 
        nc5316, nc5317, nc5318, nc5319, nc5320, nc5321, nc5322, nc5323, 
        nc5324, \A_DOUT_TEMPR110[9] , \A_DOUT_TEMPR110[8] , 
        \A_DOUT_TEMPR110[7] , \A_DOUT_TEMPR110[6] , 
        \A_DOUT_TEMPR110[5] }), .B_DOUT({nc5325, nc5326, nc5327, 
        nc5328, nc5329, nc5330, nc5331, nc5332, nc5333, nc5334, nc5335, 
        nc5336, nc5337, nc5338, nc5339, \B_DOUT_TEMPR110[9] , 
        \B_DOUT_TEMPR110[8] , \B_DOUT_TEMPR110[7] , 
        \B_DOUT_TEMPR110[6] , \B_DOUT_TEMPR110[5] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[110][1] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[9], 
        B_DIN[8], B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1818 (.A(\A_DOUT_TEMPR115[25] ), .B(\A_DOUT_TEMPR116[25] ), 
        .C(\A_DOUT_TEMPR117[25] ), .D(\A_DOUT_TEMPR118[25] ), .Y(
        OR4_1818_Y));
    OR4 OR4_417 (.A(\A_DOUT_TEMPR20[27] ), .B(\A_DOUT_TEMPR21[27] ), 
        .C(\A_DOUT_TEMPR22[27] ), .D(\A_DOUT_TEMPR23[27] ), .Y(
        OR4_417_Y));
    OR4 OR4_571 (.A(\B_DOUT_TEMPR44[9] ), .B(\B_DOUT_TEMPR45[9] ), .C(
        \B_DOUT_TEMPR46[9] ), .D(\B_DOUT_TEMPR47[9] ), .Y(OR4_571_Y));
    OR4 OR4_578 (.A(\A_DOUT_TEMPR103[5] ), .B(\A_DOUT_TEMPR104[5] ), 
        .C(\A_DOUT_TEMPR105[5] ), .D(\A_DOUT_TEMPR106[5] ), .Y(
        OR4_578_Y));
    OR4 OR4_129 (.A(\B_DOUT_TEMPR16[17] ), .B(\B_DOUT_TEMPR17[17] ), 
        .C(\B_DOUT_TEMPR18[17] ), .D(\B_DOUT_TEMPR19[17] ), .Y(
        OR4_129_Y));
    OR4 OR4_752 (.A(\B_DOUT_TEMPR12[21] ), .B(\B_DOUT_TEMPR13[21] ), 
        .C(\B_DOUT_TEMPR14[21] ), .D(\B_DOUT_TEMPR15[21] ), .Y(
        OR4_752_Y));
    OR4 OR4_356 (.A(\B_DOUT_TEMPR68[24] ), .B(\B_DOUT_TEMPR69[24] ), 
        .C(\B_DOUT_TEMPR70[24] ), .D(\B_DOUT_TEMPR71[24] ), .Y(
        OR4_356_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%90%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R90C2 (
        .A_DOUT({nc5340, nc5341, nc5342, nc5343, nc5344, nc5345, 
        nc5346, nc5347, nc5348, nc5349, nc5350, nc5351, nc5352, nc5353, 
        nc5354, \A_DOUT_TEMPR90[14] , \A_DOUT_TEMPR90[13] , 
        \A_DOUT_TEMPR90[12] , \A_DOUT_TEMPR90[11] , 
        \A_DOUT_TEMPR90[10] }), .B_DOUT({nc5355, nc5356, nc5357, 
        nc5358, nc5359, nc5360, nc5361, nc5362, nc5363, nc5364, nc5365, 
        nc5366, nc5367, nc5368, nc5369, \B_DOUT_TEMPR90[14] , 
        \B_DOUT_TEMPR90[13] , \B_DOUT_TEMPR90[12] , 
        \B_DOUT_TEMPR90[11] , \B_DOUT_TEMPR90[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[90][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2960 (.A(\B_DOUT_TEMPR44[2] ), .B(\B_DOUT_TEMPR45[2] ), .C(
        \B_DOUT_TEMPR46[2] ), .D(\B_DOUT_TEMPR47[2] ), .Y(OR4_2960_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%13%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R13C5 (
        .A_DOUT({nc5370, nc5371, nc5372, nc5373, nc5374, nc5375, 
        nc5376, nc5377, nc5378, nc5379, nc5380, nc5381, nc5382, nc5383, 
        nc5384, \A_DOUT_TEMPR13[29] , \A_DOUT_TEMPR13[28] , 
        \A_DOUT_TEMPR13[27] , \A_DOUT_TEMPR13[26] , 
        \A_DOUT_TEMPR13[25] }), .B_DOUT({nc5385, nc5386, nc5387, 
        nc5388, nc5389, nc5390, nc5391, nc5392, nc5393, nc5394, nc5395, 
        nc5396, nc5397, nc5398, nc5399, \B_DOUT_TEMPR13[29] , 
        \B_DOUT_TEMPR13[28] , \B_DOUT_TEMPR13[27] , 
        \B_DOUT_TEMPR13[26] , \B_DOUT_TEMPR13[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[13][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_706 (.A(\B_DOUT_TEMPR32[26] ), .B(\B_DOUT_TEMPR33[26] ), 
        .C(\B_DOUT_TEMPR34[26] ), .D(\B_DOUT_TEMPR35[26] ), .Y(
        OR4_706_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%8%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R8C0 (
        .A_DOUT({nc5400, nc5401, nc5402, nc5403, nc5404, nc5405, 
        nc5406, nc5407, nc5408, nc5409, nc5410, nc5411, nc5412, nc5413, 
        nc5414, \A_DOUT_TEMPR8[4] , \A_DOUT_TEMPR8[3] , 
        \A_DOUT_TEMPR8[2] , \A_DOUT_TEMPR8[1] , \A_DOUT_TEMPR8[0] }), 
        .B_DOUT({nc5415, nc5416, nc5417, nc5418, nc5419, nc5420, 
        nc5421, nc5422, nc5423, nc5424, nc5425, nc5426, nc5427, nc5428, 
        nc5429, \B_DOUT_TEMPR8[4] , \B_DOUT_TEMPR8[3] , 
        \B_DOUT_TEMPR8[2] , \B_DOUT_TEMPR8[1] , \B_DOUT_TEMPR8[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[8][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2446 (.A(\B_DOUT_TEMPR32[2] ), .B(\B_DOUT_TEMPR33[2] ), .C(
        \B_DOUT_TEMPR34[2] ), .D(\B_DOUT_TEMPR35[2] ), .Y(OR4_2446_Y));
    OR4 OR4_440 (.A(OR4_744_Y), .B(OR4_219_Y), .C(OR4_1553_Y), .D(
        OR4_2480_Y), .Y(OR4_440_Y));
    OR4 OR4_2390 (.A(\A_DOUT_TEMPR83[12] ), .B(\A_DOUT_TEMPR84[12] ), 
        .C(\A_DOUT_TEMPR85[12] ), .D(\A_DOUT_TEMPR86[12] ), .Y(
        OR4_2390_Y));
    OR4 OR4_2489 (.A(\A_DOUT_TEMPR4[7] ), .B(\A_DOUT_TEMPR5[7] ), .C(
        \A_DOUT_TEMPR6[7] ), .D(\A_DOUT_TEMPR7[7] ), .Y(OR4_2489_Y));
    OR4 OR4_557 (.A(OR4_2853_Y), .B(OR4_2144_Y), .C(OR4_1061_Y), .D(
        OR4_1067_Y), .Y(OR4_557_Y));
    OR4 OR4_2497 (.A(\B_DOUT_TEMPR36[12] ), .B(\B_DOUT_TEMPR37[12] ), 
        .C(\B_DOUT_TEMPR38[12] ), .D(\B_DOUT_TEMPR39[12] ), .Y(
        OR4_2497_Y));
    OR4 OR4_375 (.A(\A_DOUT_TEMPR95[11] ), .B(\A_DOUT_TEMPR96[11] ), 
        .C(\A_DOUT_TEMPR97[11] ), .D(\A_DOUT_TEMPR98[11] ), .Y(
        OR4_375_Y));
    OR4 OR4_1029 (.A(OR4_1722_Y), .B(OR4_2945_Y), .C(OR2_29_Y), .D(
        \B_DOUT_TEMPR74[10] ), .Y(OR4_1029_Y));
    OR4 OR4_2378 (.A(OR4_1041_Y), .B(OR4_2185_Y), .C(OR4_207_Y), .D(
        OR4_2059_Y), .Y(OR4_2378_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%78%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R78C2 (
        .A_DOUT({nc5430, nc5431, nc5432, nc5433, nc5434, nc5435, 
        nc5436, nc5437, nc5438, nc5439, nc5440, nc5441, nc5442, nc5443, 
        nc5444, \A_DOUT_TEMPR78[14] , \A_DOUT_TEMPR78[13] , 
        \A_DOUT_TEMPR78[12] , \A_DOUT_TEMPR78[11] , 
        \A_DOUT_TEMPR78[10] }), .B_DOUT({nc5445, nc5446, nc5447, 
        nc5448, nc5449, nc5450, nc5451, nc5452, nc5453, nc5454, nc5455, 
        nc5456, nc5457, nc5458, nc5459, \B_DOUT_TEMPR78[14] , 
        \B_DOUT_TEMPR78[13] , \B_DOUT_TEMPR78[12] , 
        \B_DOUT_TEMPR78[11] , \B_DOUT_TEMPR78[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[78][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1802 (.A(\A_DOUT_TEMPR115[20] ), .B(\A_DOUT_TEMPR116[20] ), 
        .C(\A_DOUT_TEMPR117[20] ), .D(\A_DOUT_TEMPR118[20] ), .Y(
        OR4_1802_Y));
    OR4 OR4_1685 (.A(\B_DOUT_TEMPR0[29] ), .B(\B_DOUT_TEMPR1[29] ), .C(
        \B_DOUT_TEMPR2[29] ), .D(\B_DOUT_TEMPR3[29] ), .Y(OR4_1685_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%68%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R68C4 (
        .A_DOUT({nc5460, nc5461, nc5462, nc5463, nc5464, nc5465, 
        nc5466, nc5467, nc5468, nc5469, nc5470, nc5471, nc5472, nc5473, 
        nc5474, \A_DOUT_TEMPR68[24] , \A_DOUT_TEMPR68[23] , 
        \A_DOUT_TEMPR68[22] , \A_DOUT_TEMPR68[21] , 
        \A_DOUT_TEMPR68[20] }), .B_DOUT({nc5475, nc5476, nc5477, 
        nc5478, nc5479, nc5480, nc5481, nc5482, nc5483, nc5484, nc5485, 
        nc5486, nc5487, nc5488, nc5489, \B_DOUT_TEMPR68[24] , 
        \B_DOUT_TEMPR68[23] , \B_DOUT_TEMPR68[22] , 
        \B_DOUT_TEMPR68[21] , \B_DOUT_TEMPR68[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[68][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_883 (.A(\A_DOUT_TEMPR32[6] ), .B(\A_DOUT_TEMPR33[6] ), .C(
        \A_DOUT_TEMPR34[6] ), .D(\A_DOUT_TEMPR35[6] ), .Y(OR4_883_Y));
    OR4 OR4_2858 (.A(\B_DOUT_TEMPR95[12] ), .B(\B_DOUT_TEMPR96[12] ), 
        .C(\B_DOUT_TEMPR97[12] ), .D(\B_DOUT_TEMPR98[12] ), .Y(
        OR4_2858_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%53%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R53C4 (
        .A_DOUT({nc5490, nc5491, nc5492, nc5493, nc5494, nc5495, 
        nc5496, nc5497, nc5498, nc5499, nc5500, nc5501, nc5502, nc5503, 
        nc5504, \A_DOUT_TEMPR53[24] , \A_DOUT_TEMPR53[23] , 
        \A_DOUT_TEMPR53[22] , \A_DOUT_TEMPR53[21] , 
        \A_DOUT_TEMPR53[20] }), .B_DOUT({nc5505, nc5506, nc5507, 
        nc5508, nc5509, nc5510, nc5511, nc5512, nc5513, nc5514, nc5515, 
        nc5516, nc5517, nc5518, nc5519, \B_DOUT_TEMPR53[24] , 
        \B_DOUT_TEMPR53[23] , \B_DOUT_TEMPR53[22] , 
        \B_DOUT_TEMPR53[21] , \B_DOUT_TEMPR53[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[53][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2762 (.A(\A_DOUT_TEMPR91[18] ), .B(\A_DOUT_TEMPR92[18] ), 
        .C(\A_DOUT_TEMPR93[18] ), .D(\A_DOUT_TEMPR94[18] ), .Y(
        OR4_2762_Y));
    OR4 OR4_1529 (.A(\B_DOUT_TEMPR56[34] ), .B(\B_DOUT_TEMPR57[34] ), 
        .C(\B_DOUT_TEMPR58[34] ), .D(\B_DOUT_TEMPR59[34] ), .Y(
        OR4_1529_Y));
    OR2 OR2_29 (.A(\B_DOUT_TEMPR72[10] ), .B(\B_DOUT_TEMPR73[10] ), .Y(
        OR2_29_Y));
    OR4 \OR4_B_DOUT[13]  (.A(OR4_1096_Y), .B(OR4_792_Y), .C(OR4_2942_Y)
        , .D(OR4_493_Y), .Y(B_DOUT[13]));
    OR4 OR4_2745 (.A(\B_DOUT_TEMPR111[36] ), .B(\B_DOUT_TEMPR112[36] ), 
        .C(\B_DOUT_TEMPR113[36] ), .D(\B_DOUT_TEMPR114[36] ), .Y(
        OR4_2745_Y));
    OR4 OR4_1194 (.A(\A_DOUT_TEMPR107[39] ), .B(\A_DOUT_TEMPR108[39] ), 
        .C(\A_DOUT_TEMPR109[39] ), .D(\A_DOUT_TEMPR110[39] ), .Y(
        OR4_1194_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%16%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R16C4 (
        .A_DOUT({nc5520, nc5521, nc5522, nc5523, nc5524, nc5525, 
        nc5526, nc5527, nc5528, nc5529, nc5530, nc5531, nc5532, nc5533, 
        nc5534, \A_DOUT_TEMPR16[24] , \A_DOUT_TEMPR16[23] , 
        \A_DOUT_TEMPR16[22] , \A_DOUT_TEMPR16[21] , 
        \A_DOUT_TEMPR16[20] }), .B_DOUT({nc5535, nc5536, nc5537, 
        nc5538, nc5539, nc5540, nc5541, nc5542, nc5543, nc5544, nc5545, 
        nc5546, nc5547, nc5548, nc5549, \B_DOUT_TEMPR16[24] , 
        \B_DOUT_TEMPR16[23] , \B_DOUT_TEMPR16[22] , 
        \B_DOUT_TEMPR16[21] , \B_DOUT_TEMPR16[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[16][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2380 (.A(\A_DOUT_TEMPR56[13] ), .B(\A_DOUT_TEMPR57[13] ), 
        .C(\A_DOUT_TEMPR58[13] ), .D(\A_DOUT_TEMPR59[13] ), .Y(
        OR4_2380_Y));
    OR4 OR4_501 (.A(OR4_1640_Y), .B(OR4_808_Y), .C(OR4_1440_Y), .D(
        OR4_631_Y), .Y(OR4_501_Y));
    OR4 OR4_2487 (.A(OR4_1233_Y), .B(OR4_2391_Y), .C(OR4_406_Y), .D(
        OR4_1811_Y), .Y(OR4_2487_Y));
    OR4 OR4_508 (.A(\B_DOUT_TEMPR20[25] ), .B(\B_DOUT_TEMPR21[25] ), 
        .C(\B_DOUT_TEMPR22[25] ), .D(\B_DOUT_TEMPR23[25] ), .Y(
        OR4_508_Y));
    OR4 OR4_1358 (.A(\B_DOUT_TEMPR52[35] ), .B(\B_DOUT_TEMPR53[35] ), 
        .C(\B_DOUT_TEMPR54[35] ), .D(\B_DOUT_TEMPR55[35] ), .Y(
        OR4_1358_Y));
    OR4 OR4_1718 (.A(OR4_1074_Y), .B(OR4_2220_Y), .C(OR4_242_Y), .D(
        OR4_2966_Y), .Y(OR4_1718_Y));
    OR4 OR4_1322 (.A(OR4_2065_Y), .B(OR4_523_Y), .C(OR4_1114_Y), .D(
        OR4_931_Y), .Y(OR4_1322_Y));
    OR4 OR4_721 (.A(OR4_193_Y), .B(OR4_2241_Y), .C(OR4_2461_Y), .D(
        OR4_2257_Y), .Y(OR4_721_Y));
    OR2 OR2_43 (.A(\B_DOUT_TEMPR72[23] ), .B(\B_DOUT_TEMPR73[23] ), .Y(
        OR2_43_Y));
    OR4 \OR4_B_DOUT[30]  (.A(OR4_105_Y), .B(OR4_2593_Y), .C(OR4_2277_Y)
        , .D(OR4_748_Y), .Y(B_DOUT[30]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%78%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R78C3 (
        .A_DOUT({nc5550, nc5551, nc5552, nc5553, nc5554, nc5555, 
        nc5556, nc5557, nc5558, nc5559, nc5560, nc5561, nc5562, nc5563, 
        nc5564, \A_DOUT_TEMPR78[19] , \A_DOUT_TEMPR78[18] , 
        \A_DOUT_TEMPR78[17] , \A_DOUT_TEMPR78[16] , 
        \A_DOUT_TEMPR78[15] }), .B_DOUT({nc5565, nc5566, nc5567, 
        nc5568, nc5569, nc5570, nc5571, nc5572, nc5573, nc5574, nc5575, 
        nc5576, nc5577, nc5578, nc5579, \B_DOUT_TEMPR78[19] , 
        \B_DOUT_TEMPR78[18] , \B_DOUT_TEMPR78[17] , 
        \B_DOUT_TEMPR78[16] , \B_DOUT_TEMPR78[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[78][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1687 (.A(OR4_578_Y), .B(OR4_2004_Y), .C(OR4_1488_Y), .D(
        OR4_2971_Y), .Y(OR4_1687_Y));
    OR4 OR4_293 (.A(\A_DOUT_TEMPR83[36] ), .B(\A_DOUT_TEMPR84[36] ), 
        .C(\A_DOUT_TEMPR85[36] ), .D(\A_DOUT_TEMPR86[36] ), .Y(
        OR4_293_Y));
    OR4 OR4_2662 (.A(\B_DOUT_TEMPR95[34] ), .B(\B_DOUT_TEMPR96[34] ), 
        .C(\B_DOUT_TEMPR97[34] ), .D(\B_DOUT_TEMPR98[34] ), .Y(
        OR4_2662_Y));
    OR4 OR4_2230 (.A(\B_DOUT_TEMPR115[30] ), .B(\B_DOUT_TEMPR116[30] ), 
        .C(\B_DOUT_TEMPR117[30] ), .D(\B_DOUT_TEMPR118[30] ), .Y(
        OR4_2230_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%15%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R15C5 (
        .A_DOUT({nc5580, nc5581, nc5582, nc5583, nc5584, nc5585, 
        nc5586, nc5587, nc5588, nc5589, nc5590, nc5591, nc5592, nc5593, 
        nc5594, \A_DOUT_TEMPR15[29] , \A_DOUT_TEMPR15[28] , 
        \A_DOUT_TEMPR15[27] , \A_DOUT_TEMPR15[26] , 
        \A_DOUT_TEMPR15[25] }), .B_DOUT({nc5595, nc5596, nc5597, 
        nc5598, nc5599, nc5600, nc5601, nc5602, nc5603, nc5604, nc5605, 
        nc5606, nc5607, nc5608, nc5609, \B_DOUT_TEMPR15[29] , 
        \B_DOUT_TEMPR15[28] , \B_DOUT_TEMPR15[27] , 
        \B_DOUT_TEMPR15[26] , \B_DOUT_TEMPR15[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[15][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1479 (.A(\B_DOUT_TEMPR95[29] ), .B(\B_DOUT_TEMPR96[29] ), 
        .C(\B_DOUT_TEMPR97[29] ), .D(\B_DOUT_TEMPR98[29] ), .Y(
        OR4_1479_Y));
    OR4 OR4_1603 (.A(OR4_153_Y), .B(OR4_920_Y), .C(OR4_443_Y), .D(
        OR4_2418_Y), .Y(OR4_1603_Y));
    OR4 OR4_182 (.A(OR4_2910_Y), .B(OR4_1511_Y), .C(OR4_905_Y), .D(
        OR4_209_Y), .Y(OR4_182_Y));
    OR4 OR4_391 (.A(\B_DOUT_TEMPR20[12] ), .B(\B_DOUT_TEMPR21[12] ), 
        .C(\B_DOUT_TEMPR22[12] ), .D(\B_DOUT_TEMPR23[12] ), .Y(
        OR4_391_Y));
    OR4 OR4_870 (.A(OR4_1314_Y), .B(OR4_2749_Y), .C(OR4_2193_Y), .D(
        OR4_246_Y), .Y(OR4_870_Y));
    OR4 OR4_895 (.A(\B_DOUT_TEMPR40[20] ), .B(\B_DOUT_TEMPR41[20] ), 
        .C(\B_DOUT_TEMPR42[20] ), .D(\B_DOUT_TEMPR43[20] ), .Y(
        OR4_895_Y));
    OR4 OR4_149 (.A(\B_DOUT_TEMPR16[2] ), .B(\B_DOUT_TEMPR17[2] ), .C(
        \B_DOUT_TEMPR18[2] ), .D(\B_DOUT_TEMPR19[2] ), .Y(OR4_149_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%74%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R74C1 (
        .A_DOUT({nc5610, nc5611, nc5612, nc5613, nc5614, nc5615, 
        nc5616, nc5617, nc5618, nc5619, nc5620, nc5621, nc5622, nc5623, 
        nc5624, \A_DOUT_TEMPR74[9] , \A_DOUT_TEMPR74[8] , 
        \A_DOUT_TEMPR74[7] , \A_DOUT_TEMPR74[6] , \A_DOUT_TEMPR74[5] })
        , .B_DOUT({nc5625, nc5626, nc5627, nc5628, nc5629, nc5630, 
        nc5631, nc5632, nc5633, nc5634, nc5635, nc5636, nc5637, nc5638, 
        nc5639, \B_DOUT_TEMPR74[9] , \B_DOUT_TEMPR74[8] , 
        \B_DOUT_TEMPR74[7] , \B_DOUT_TEMPR74[6] , \B_DOUT_TEMPR74[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[74][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%14%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R14C5 (
        .A_DOUT({nc5640, nc5641, nc5642, nc5643, nc5644, nc5645, 
        nc5646, nc5647, nc5648, nc5649, nc5650, nc5651, nc5652, nc5653, 
        nc5654, \A_DOUT_TEMPR14[29] , \A_DOUT_TEMPR14[28] , 
        \A_DOUT_TEMPR14[27] , \A_DOUT_TEMPR14[26] , 
        \A_DOUT_TEMPR14[25] }), .B_DOUT({nc5655, nc5656, nc5657, 
        nc5658, nc5659, nc5660, nc5661, nc5662, nc5663, nc5664, nc5665, 
        nc5666, nc5667, nc5668, nc5669, \B_DOUT_TEMPR14[29] , 
        \B_DOUT_TEMPR14[28] , \B_DOUT_TEMPR14[27] , 
        \B_DOUT_TEMPR14[26] , \B_DOUT_TEMPR14[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[14][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1909 (.A(OR4_533_Y), .B(OR4_48_Y), .C(OR4_2236_Y), .D(
        OR4_1211_Y), .Y(OR4_1909_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%70%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R70C4 (
        .A_DOUT({nc5670, nc5671, nc5672, nc5673, nc5674, nc5675, 
        nc5676, nc5677, nc5678, nc5679, nc5680, nc5681, nc5682, nc5683, 
        nc5684, \A_DOUT_TEMPR70[24] , \A_DOUT_TEMPR70[23] , 
        \A_DOUT_TEMPR70[22] , \A_DOUT_TEMPR70[21] , 
        \A_DOUT_TEMPR70[20] }), .B_DOUT({nc5685, nc5686, nc5687, 
        nc5688, nc5689, nc5690, nc5691, nc5692, nc5693, nc5694, nc5695, 
        nc5696, nc5697, nc5698, nc5699, \B_DOUT_TEMPR70[24] , 
        \B_DOUT_TEMPR70[23] , \B_DOUT_TEMPR70[22] , 
        \B_DOUT_TEMPR70[21] , \B_DOUT_TEMPR70[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[70][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_193 (.A(\B_DOUT_TEMPR48[16] ), .B(\B_DOUT_TEMPR49[16] ), 
        .C(\B_DOUT_TEMPR50[16] ), .D(\B_DOUT_TEMPR51[16] ), .Y(
        OR4_193_Y));
    OR4 OR4_1230 (.A(\B_DOUT_TEMPR91[21] ), .B(\B_DOUT_TEMPR92[21] ), 
        .C(\B_DOUT_TEMPR93[21] ), .D(\B_DOUT_TEMPR94[21] ), .Y(
        OR4_1230_Y));
    OR4 OR4_570 (.A(OR4_152_Y), .B(OR4_412_Y), .C(OR4_1891_Y), .D(
        OR4_414_Y), .Y(OR4_570_Y));
    OR4 OR4_2962 (.A(\B_DOUT_TEMPR8[31] ), .B(\B_DOUT_TEMPR9[31] ), .C(
        \B_DOUT_TEMPR10[31] ), .D(\B_DOUT_TEMPR11[31] ), .Y(OR4_2962_Y)
        );
    OR2 OR2_62 (.A(\B_DOUT_TEMPR72[2] ), .B(\B_DOUT_TEMPR73[2] ), .Y(
        OR2_62_Y));
    OR4 OR4_2625 (.A(\A_DOUT_TEMPR36[11] ), .B(\A_DOUT_TEMPR37[11] ), 
        .C(\A_DOUT_TEMPR38[11] ), .D(\A_DOUT_TEMPR39[11] ), .Y(
        OR4_2625_Y));
    OR4 OR4_1895 (.A(\A_DOUT_TEMPR20[16] ), .B(\A_DOUT_TEMPR21[16] ), 
        .C(\A_DOUT_TEMPR22[16] ), .D(\A_DOUT_TEMPR23[16] ), .Y(
        OR4_1895_Y));
    OR4 OR4_305 (.A(\B_DOUT_TEMPR87[36] ), .B(\B_DOUT_TEMPR88[36] ), 
        .C(\B_DOUT_TEMPR89[36] ), .D(\B_DOUT_TEMPR90[36] ), .Y(
        OR4_305_Y));
    OR4 OR4_985 (.A(\B_DOUT_TEMPR40[2] ), .B(\B_DOUT_TEMPR41[2] ), .C(
        \B_DOUT_TEMPR42[2] ), .D(\B_DOUT_TEMPR43[2] ), .Y(OR4_985_Y));
    OR4 OR4_485 (.A(\B_DOUT_TEMPR91[27] ), .B(\B_DOUT_TEMPR92[27] ), 
        .C(\B_DOUT_TEMPR93[27] ), .D(\B_DOUT_TEMPR94[27] ), .Y(
        OR4_485_Y));
    OR4 OR4_822 (.A(\B_DOUT_TEMPR8[5] ), .B(\B_DOUT_TEMPR9[5] ), .C(
        \B_DOUT_TEMPR10[5] ), .D(\B_DOUT_TEMPR11[5] ), .Y(OR4_822_Y));
    OR4 OR4_2475 (.A(\A_DOUT_TEMPR28[20] ), .B(\A_DOUT_TEMPR29[20] ), 
        .C(\A_DOUT_TEMPR30[20] ), .D(\A_DOUT_TEMPR31[20] ), .Y(
        OR4_2475_Y));
    OR2 OR2_12 (.A(\B_DOUT_TEMPR72[14] ), .B(\B_DOUT_TEMPR73[14] ), .Y(
        OR2_12_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%51%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R51C4 (
        .A_DOUT({nc5700, nc5701, nc5702, nc5703, nc5704, nc5705, 
        nc5706, nc5707, nc5708, nc5709, nc5710, nc5711, nc5712, nc5713, 
        nc5714, \A_DOUT_TEMPR51[24] , \A_DOUT_TEMPR51[23] , 
        \A_DOUT_TEMPR51[22] , \A_DOUT_TEMPR51[21] , 
        \A_DOUT_TEMPR51[20] }), .B_DOUT({nc5715, nc5716, nc5717, 
        nc5718, nc5719, nc5720, nc5721, nc5722, nc5723, nc5724, nc5725, 
        nc5726, nc5727, nc5728, nc5729, \B_DOUT_TEMPR51[24] , 
        \B_DOUT_TEMPR51[23] , \B_DOUT_TEMPR51[22] , 
        \B_DOUT_TEMPR51[21] , \B_DOUT_TEMPR51[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[51][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2758 (.A(\A_DOUT_TEMPR56[8] ), .B(\A_DOUT_TEMPR57[8] ), .C(
        \A_DOUT_TEMPR58[8] ), .D(\A_DOUT_TEMPR59[8] ), .Y(OR4_2758_Y));
    OR4 OR4_774 (.A(\A_DOUT_TEMPR48[20] ), .B(\A_DOUT_TEMPR49[20] ), 
        .C(\A_DOUT_TEMPR50[20] ), .D(\A_DOUT_TEMPR51[20] ), .Y(
        OR4_774_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%105%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R105C0 (
        .A_DOUT({nc5730, nc5731, nc5732, nc5733, nc5734, nc5735, 
        nc5736, nc5737, nc5738, nc5739, nc5740, nc5741, nc5742, nc5743, 
        nc5744, \A_DOUT_TEMPR105[4] , \A_DOUT_TEMPR105[3] , 
        \A_DOUT_TEMPR105[2] , \A_DOUT_TEMPR105[1] , 
        \A_DOUT_TEMPR105[0] }), .B_DOUT({nc5745, nc5746, nc5747, 
        nc5748, nc5749, nc5750, nc5751, nc5752, nc5753, nc5754, nc5755, 
        nc5756, nc5757, nc5758, nc5759, \B_DOUT_TEMPR105[4] , 
        \B_DOUT_TEMPR105[3] , \B_DOUT_TEMPR105[2] , 
        \B_DOUT_TEMPR105[1] , \B_DOUT_TEMPR105[0] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[105][0] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[4], 
        B_DIN[3], B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1525 (.A(OR4_186_Y), .B(OR4_1682_Y), .C(OR4_2251_Y), .D(
        OR4_2083_Y), .Y(OR4_1525_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%106%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R106C4 (
        .A_DOUT({nc5760, nc5761, nc5762, nc5763, nc5764, nc5765, 
        nc5766, nc5767, nc5768, nc5769, nc5770, nc5771, nc5772, nc5773, 
        nc5774, \A_DOUT_TEMPR106[24] , \A_DOUT_TEMPR106[23] , 
        \A_DOUT_TEMPR106[22] , \A_DOUT_TEMPR106[21] , 
        \A_DOUT_TEMPR106[20] }), .B_DOUT({nc5775, nc5776, nc5777, 
        nc5778, nc5779, nc5780, nc5781, nc5782, nc5783, nc5784, nc5785, 
        nc5786, nc5787, nc5788, nc5789, \B_DOUT_TEMPR106[24] , 
        \B_DOUT_TEMPR106[23] , \B_DOUT_TEMPR106[22] , 
        \B_DOUT_TEMPR106[21] , \B_DOUT_TEMPR106[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[106][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2336 (.A(\B_DOUT_TEMPR8[9] ), .B(\B_DOUT_TEMPR9[9] ), .C(
        \B_DOUT_TEMPR10[9] ), .D(\B_DOUT_TEMPR11[9] ), .Y(OR4_2336_Y));
    OR4 OR4_1848 (.A(\B_DOUT_TEMPR60[2] ), .B(\B_DOUT_TEMPR61[2] ), .C(
        \B_DOUT_TEMPR62[2] ), .D(\B_DOUT_TEMPR63[2] ), .Y(OR4_1848_Y));
    OR4 OR4_1370 (.A(\A_DOUT_TEMPR36[0] ), .B(\A_DOUT_TEMPR37[0] ), .C(
        \A_DOUT_TEMPR38[0] ), .D(\A_DOUT_TEMPR39[0] ), .Y(OR4_1370_Y));
    OR4 OR4_2108 (.A(\A_DOUT_TEMPR103[3] ), .B(\A_DOUT_TEMPR104[3] ), 
        .C(\A_DOUT_TEMPR105[3] ), .D(\A_DOUT_TEMPR106[3] ), .Y(
        OR4_2108_Y));
    OR4 OR4_1477 (.A(\B_DOUT_TEMPR95[0] ), .B(\B_DOUT_TEMPR96[0] ), .C(
        \B_DOUT_TEMPR97[0] ), .D(\B_DOUT_TEMPR98[0] ), .Y(OR4_1477_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%64%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R64C7 (
        .A_DOUT({nc5790, nc5791, nc5792, nc5793, nc5794, nc5795, 
        nc5796, nc5797, nc5798, nc5799, nc5800, nc5801, nc5802, nc5803, 
        nc5804, \A_DOUT_TEMPR64[39] , \A_DOUT_TEMPR64[38] , 
        \A_DOUT_TEMPR64[37] , \A_DOUT_TEMPR64[36] , 
        \A_DOUT_TEMPR64[35] }), .B_DOUT({nc5805, nc5806, nc5807, 
        nc5808, nc5809, nc5810, nc5811, nc5812, nc5813, nc5814, nc5815, 
        nc5816, nc5817, nc5818, nc5819, \B_DOUT_TEMPR64[39] , 
        \B_DOUT_TEMPR64[38] , \B_DOUT_TEMPR64[37] , 
        \B_DOUT_TEMPR64[36] , \B_DOUT_TEMPR64[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[64][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%33%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R33C4 (
        .A_DOUT({nc5820, nc5821, nc5822, nc5823, nc5824, nc5825, 
        nc5826, nc5827, nc5828, nc5829, nc5830, nc5831, nc5832, nc5833, 
        nc5834, \A_DOUT_TEMPR33[24] , \A_DOUT_TEMPR33[23] , 
        \A_DOUT_TEMPR33[22] , \A_DOUT_TEMPR33[21] , 
        \A_DOUT_TEMPR33[20] }), .B_DOUT({nc5835, nc5836, nc5837, 
        nc5838, nc5839, nc5840, nc5841, nc5842, nc5843, nc5844, nc5845, 
        nc5846, nc5847, nc5848, nc5849, \B_DOUT_TEMPR33[24] , 
        \B_DOUT_TEMPR33[23] , \B_DOUT_TEMPR33[22] , 
        \B_DOUT_TEMPR33[21] , \B_DOUT_TEMPR33[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[33][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%117%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R117C7 (
        .A_DOUT({nc5850, nc5851, nc5852, nc5853, nc5854, nc5855, 
        nc5856, nc5857, nc5858, nc5859, nc5860, nc5861, nc5862, nc5863, 
        nc5864, \A_DOUT_TEMPR117[39] , \A_DOUT_TEMPR117[38] , 
        \A_DOUT_TEMPR117[37] , \A_DOUT_TEMPR117[36] , 
        \A_DOUT_TEMPR117[35] }), .B_DOUT({nc5865, nc5866, nc5867, 
        nc5868, nc5869, nc5870, nc5871, nc5872, nc5873, nc5874, nc5875, 
        nc5876, nc5877, nc5878, nc5879, \B_DOUT_TEMPR117[39] , 
        \B_DOUT_TEMPR117[38] , \B_DOUT_TEMPR117[37] , 
        \B_DOUT_TEMPR117[36] , \B_DOUT_TEMPR117[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[117][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1704 (.A(\A_DOUT_TEMPR91[30] ), .B(\A_DOUT_TEMPR92[30] ), 
        .C(\A_DOUT_TEMPR93[30] ), .D(\A_DOUT_TEMPR94[30] ), .Y(
        OR4_1704_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%41%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R41C2 (
        .A_DOUT({nc5880, nc5881, nc5882, nc5883, nc5884, nc5885, 
        nc5886, nc5887, nc5888, nc5889, nc5890, nc5891, nc5892, nc5893, 
        nc5894, \A_DOUT_TEMPR41[14] , \A_DOUT_TEMPR41[13] , 
        \A_DOUT_TEMPR41[12] , \A_DOUT_TEMPR41[11] , 
        \A_DOUT_TEMPR41[10] }), .B_DOUT({nc5895, nc5896, nc5897, 
        nc5898, nc5899, nc5900, nc5901, nc5902, nc5903, nc5904, nc5905, 
        nc5906, nc5907, nc5908, nc5909, \B_DOUT_TEMPR41[14] , 
        \B_DOUT_TEMPR41[13] , \B_DOUT_TEMPR41[12] , 
        \B_DOUT_TEMPR41[11] , \B_DOUT_TEMPR41[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[41][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1336 (.A(\B_DOUT_TEMPR24[14] ), .B(\B_DOUT_TEMPR25[14] ), 
        .C(\B_DOUT_TEMPR26[14] ), .D(\B_DOUT_TEMPR27[14] ), .Y(
        OR4_1336_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%94%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R94C6 (
        .A_DOUT({nc5910, nc5911, nc5912, nc5913, nc5914, nc5915, 
        nc5916, nc5917, nc5918, nc5919, nc5920, nc5921, nc5922, nc5923, 
        nc5924, \A_DOUT_TEMPR94[34] , \A_DOUT_TEMPR94[33] , 
        \A_DOUT_TEMPR94[32] , \A_DOUT_TEMPR94[31] , 
        \A_DOUT_TEMPR94[30] }), .B_DOUT({nc5925, nc5926, nc5927, 
        nc5928, nc5929, nc5930, nc5931, nc5932, nc5933, nc5934, nc5935, 
        nc5936, nc5937, nc5938, nc5939, \B_DOUT_TEMPR94[34] , 
        \B_DOUT_TEMPR94[33] , \B_DOUT_TEMPR94[32] , 
        \B_DOUT_TEMPR94[31] , \B_DOUT_TEMPR94[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[94][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1562 (.A(\B_DOUT_TEMPR75[14] ), .B(\B_DOUT_TEMPR76[14] ), 
        .C(\B_DOUT_TEMPR77[14] ), .D(\B_DOUT_TEMPR78[14] ), .Y(
        OR4_1562_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%80%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R80C0 (
        .A_DOUT({nc5940, nc5941, nc5942, nc5943, nc5944, nc5945, 
        nc5946, nc5947, nc5948, nc5949, nc5950, nc5951, nc5952, nc5953, 
        nc5954, \A_DOUT_TEMPR80[4] , \A_DOUT_TEMPR80[3] , 
        \A_DOUT_TEMPR80[2] , \A_DOUT_TEMPR80[1] , \A_DOUT_TEMPR80[0] })
        , .B_DOUT({nc5955, nc5956, nc5957, nc5958, nc5959, nc5960, 
        nc5961, nc5962, nc5963, nc5964, nc5965, nc5966, nc5967, nc5968, 
        nc5969, \B_DOUT_TEMPR80[4] , \B_DOUT_TEMPR80[3] , 
        \B_DOUT_TEMPR80[2] , \B_DOUT_TEMPR80[1] , \B_DOUT_TEMPR80[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[80][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2627 (.A(\B_DOUT_TEMPR95[18] ), .B(\B_DOUT_TEMPR96[18] ), 
        .C(\B_DOUT_TEMPR97[18] ), .D(\B_DOUT_TEMPR98[18] ), .Y(
        OR4_2627_Y));
    OR4 OR4_792 (.A(OR4_49_Y), .B(OR4_929_Y), .C(OR4_2376_Y), .D(
        OR4_932_Y), .Y(OR4_792_Y));
    OR4 OR4_1401 (.A(\B_DOUT_TEMPR79[32] ), .B(\B_DOUT_TEMPR80[32] ), 
        .C(\B_DOUT_TEMPR81[32] ), .D(\B_DOUT_TEMPR82[32] ), .Y(
        OR4_1401_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%103%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R103C3 (
        .A_DOUT({nc5970, nc5971, nc5972, nc5973, nc5974, nc5975, 
        nc5976, nc5977, nc5978, nc5979, nc5980, nc5981, nc5982, nc5983, 
        nc5984, \A_DOUT_TEMPR103[19] , \A_DOUT_TEMPR103[18] , 
        \A_DOUT_TEMPR103[17] , \A_DOUT_TEMPR103[16] , 
        \A_DOUT_TEMPR103[15] }), .B_DOUT({nc5985, nc5986, nc5987, 
        nc5988, nc5989, nc5990, nc5991, nc5992, nc5993, nc5994, nc5995, 
        nc5996, nc5997, nc5998, nc5999, \B_DOUT_TEMPR103[19] , 
        \B_DOUT_TEMPR103[18] , \B_DOUT_TEMPR103[17] , 
        \B_DOUT_TEMPR103[16] , \B_DOUT_TEMPR103[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[103][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%85%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R85C4 (
        .A_DOUT({nc6000, nc6001, nc6002, nc6003, nc6004, nc6005, 
        nc6006, nc6007, nc6008, nc6009, nc6010, nc6011, nc6012, nc6013, 
        nc6014, \A_DOUT_TEMPR85[24] , \A_DOUT_TEMPR85[23] , 
        \A_DOUT_TEMPR85[22] , \A_DOUT_TEMPR85[21] , 
        \A_DOUT_TEMPR85[20] }), .B_DOUT({nc6015, nc6016, nc6017, 
        nc6018, nc6019, nc6020, nc6021, nc6022, nc6023, nc6024, nc6025, 
        nc6026, nc6027, nc6028, nc6029, \B_DOUT_TEMPR85[24] , 
        \B_DOUT_TEMPR85[23] , \B_DOUT_TEMPR85[22] , 
        \B_DOUT_TEMPR85[21] , \B_DOUT_TEMPR85[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[85][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_756 (.A(\B_DOUT_TEMPR75[36] ), .B(\B_DOUT_TEMPR76[36] ), 
        .C(\B_DOUT_TEMPR77[36] ), .D(\B_DOUT_TEMPR78[36] ), .Y(
        OR4_756_Y));
    OR4 OR4_1455 (.A(\B_DOUT_TEMPR64[11] ), .B(\B_DOUT_TEMPR65[11] ), 
        .C(\B_DOUT_TEMPR66[11] ), .D(\B_DOUT_TEMPR67[11] ), .Y(
        OR4_1455_Y));
    OR4 OR4_396 (.A(OR4_2395_Y), .B(OR4_1615_Y), .C(OR4_62_Y), .D(
        OR4_1616_Y), .Y(OR4_396_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%51%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R51C3 (
        .A_DOUT({nc6030, nc6031, nc6032, nc6033, nc6034, nc6035, 
        nc6036, nc6037, nc6038, nc6039, nc6040, nc6041, nc6042, nc6043, 
        nc6044, \A_DOUT_TEMPR51[19] , \A_DOUT_TEMPR51[18] , 
        \A_DOUT_TEMPR51[17] , \A_DOUT_TEMPR51[16] , 
        \A_DOUT_TEMPR51[15] }), .B_DOUT({nc6045, nc6046, nc6047, 
        nc6048, nc6049, nc6050, nc6051, nc6052, nc6053, nc6054, nc6055, 
        nc6056, nc6057, nc6058, nc6059, \B_DOUT_TEMPR51[19] , 
        \B_DOUT_TEMPR51[18] , \B_DOUT_TEMPR51[17] , 
        \B_DOUT_TEMPR51[16] , \B_DOUT_TEMPR51[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[51][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2803 (.A(\B_DOUT_TEMPR60[37] ), .B(\B_DOUT_TEMPR61[37] ), 
        .C(\B_DOUT_TEMPR62[37] ), .D(\B_DOUT_TEMPR63[37] ), .Y(
        OR4_2803_Y));
    OR4 OR4_2776 (.A(\B_DOUT_TEMPR87[15] ), .B(\B_DOUT_TEMPR88[15] ), 
        .C(\B_DOUT_TEMPR89[15] ), .D(\B_DOUT_TEMPR90[15] ), .Y(
        OR4_2776_Y));
    OR4 OR4_977 (.A(OR4_1368_Y), .B(OR4_1643_Y), .C(OR4_1304_Y), .D(
        OR4_1667_Y), .Y(OR4_977_Y));
    OR4 OR4_800 (.A(OR4_619_Y), .B(OR4_1940_Y), .C(OR4_1580_Y), .D(
        OR4_2646_Y), .Y(OR4_800_Y));
    OR4 OR4_2711 (.A(\B_DOUT_TEMPR68[33] ), .B(\B_DOUT_TEMPR69[33] ), 
        .C(\B_DOUT_TEMPR70[33] ), .D(\B_DOUT_TEMPR71[33] ), .Y(
        OR4_2711_Y));
    OR4 OR4_467 (.A(\B_DOUT_TEMPR44[19] ), .B(\B_DOUT_TEMPR45[19] ), 
        .C(\B_DOUT_TEMPR46[19] ), .D(\B_DOUT_TEMPR47[19] ), .Y(
        OR4_467_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_2 (.A(B_ADDR[16]), .B(B_ADDR[15]), .C(
        B_ADDR[14]), .Y(CFG3_2_Y));
    OR4 OR4_741 (.A(\B_DOUT_TEMPR20[3] ), .B(\B_DOUT_TEMPR21[3] ), .C(
        \B_DOUT_TEMPR22[3] ), .D(\B_DOUT_TEMPR23[3] ), .Y(OR4_741_Y));
    OR4 OR4_597 (.A(\A_DOUT_TEMPR8[5] ), .B(\A_DOUT_TEMPR9[5] ), .C(
        \A_DOUT_TEMPR10[5] ), .D(\A_DOUT_TEMPR11[5] ), .Y(OR4_597_Y));
    OR4 OR4_1384 (.A(OR4_934_Y), .B(OR4_716_Y), .C(OR2_21_Y), .D(
        \A_DOUT_TEMPR74[36] ), .Y(OR4_1384_Y));
    OR4 OR4_500 (.A(\B_DOUT_TEMPR20[13] ), .B(\B_DOUT_TEMPR21[13] ), 
        .C(\B_DOUT_TEMPR22[13] ), .D(\B_DOUT_TEMPR23[13] ), .Y(
        OR4_500_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%25%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R25C2 (
        .A_DOUT({nc6060, nc6061, nc6062, nc6063, nc6064, nc6065, 
        nc6066, nc6067, nc6068, nc6069, nc6070, nc6071, nc6072, nc6073, 
        nc6074, \A_DOUT_TEMPR25[14] , \A_DOUT_TEMPR25[13] , 
        \A_DOUT_TEMPR25[12] , \A_DOUT_TEMPR25[11] , 
        \A_DOUT_TEMPR25[10] }), .B_DOUT({nc6075, nc6076, nc6077, 
        nc6078, nc6079, nc6080, nc6081, nc6082, nc6083, nc6084, nc6085, 
        nc6086, nc6087, nc6088, nc6089, \B_DOUT_TEMPR25[14] , 
        \B_DOUT_TEMPR25[13] , \B_DOUT_TEMPR25[12] , 
        \B_DOUT_TEMPR25[11] , \B_DOUT_TEMPR25[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[25][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2709 (.A(\A_DOUT_TEMPR24[30] ), .B(\A_DOUT_TEMPR25[30] ), 
        .C(\A_DOUT_TEMPR26[30] ), .D(\A_DOUT_TEMPR27[30] ), .Y(
        OR4_2709_Y));
    OR4 OR4_2546 (.A(\B_DOUT_TEMPR44[24] ), .B(\B_DOUT_TEMPR45[24] ), 
        .C(\B_DOUT_TEMPR46[24] ), .D(\B_DOUT_TEMPR47[24] ), .Y(
        OR4_2546_Y));
    OR4 OR4_1928 (.A(OR4_1123_Y), .B(OR4_1484_Y), .C(OR4_2207_Y), .D(
        OR4_27_Y), .Y(OR4_1928_Y));
    OR4 OR4_576 (.A(OR4_2382_Y), .B(OR4_938_Y), .C(OR4_1735_Y), .D(
        OR4_764_Y), .Y(OR4_576_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%103%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R103C5 (
        .A_DOUT({nc6090, nc6091, nc6092, nc6093, nc6094, nc6095, 
        nc6096, nc6097, nc6098, nc6099, nc6100, nc6101, nc6102, nc6103, 
        nc6104, \A_DOUT_TEMPR103[29] , \A_DOUT_TEMPR103[28] , 
        \A_DOUT_TEMPR103[27] , \A_DOUT_TEMPR103[26] , 
        \A_DOUT_TEMPR103[25] }), .B_DOUT({nc6105, nc6106, nc6107, 
        nc6108, nc6109, nc6110, nc6111, nc6112, nc6113, nc6114, nc6115, 
        nc6116, nc6117, nc6118, nc6119, \B_DOUT_TEMPR103[29] , 
        \B_DOUT_TEMPR103[28] , \B_DOUT_TEMPR103[27] , 
        \B_DOUT_TEMPR103[26] , \B_DOUT_TEMPR103[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[103][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2747 (.A(\A_DOUT_TEMPR36[6] ), .B(\A_DOUT_TEMPR37[6] ), .C(
        \A_DOUT_TEMPR38[6] ), .D(\A_DOUT_TEMPR39[6] ), .Y(OR4_2747_Y));
    OR4 OR4_1756 (.A(\B_DOUT_TEMPR111[1] ), .B(\B_DOUT_TEMPR112[1] ), 
        .C(\B_DOUT_TEMPR113[1] ), .D(\B_DOUT_TEMPR114[1] ), .Y(
        OR4_1756_Y));
    OR4 OR4_704 (.A(OR4_2454_Y), .B(OR4_2790_Y), .C(OR4_2384_Y), .D(
        OR4_2805_Y), .Y(OR4_704_Y));
    OR4 OR4_2541 (.A(\B_DOUT_TEMPR32[22] ), .B(\B_DOUT_TEMPR33[22] ), 
        .C(\B_DOUT_TEMPR34[22] ), .D(\B_DOUT_TEMPR35[22] ), .Y(
        OR4_2541_Y));
    OR4 OR4_551 (.A(\B_DOUT_TEMPR48[13] ), .B(\B_DOUT_TEMPR49[13] ), 
        .C(\B_DOUT_TEMPR50[13] ), .D(\B_DOUT_TEMPR51[13] ), .Y(
        OR4_551_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%72%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R72C2 (
        .A_DOUT({nc6120, nc6121, nc6122, nc6123, nc6124, nc6125, 
        nc6126, nc6127, nc6128, nc6129, nc6130, nc6131, nc6132, nc6133, 
        nc6134, \A_DOUT_TEMPR72[14] , \A_DOUT_TEMPR72[13] , 
        \A_DOUT_TEMPR72[12] , \A_DOUT_TEMPR72[11] , 
        \A_DOUT_TEMPR72[10] }), .B_DOUT({nc6135, nc6136, nc6137, 
        nc6138, nc6139, nc6140, nc6141, nc6142, nc6143, nc6144, nc6145, 
        nc6146, nc6147, nc6148, nc6149, \B_DOUT_TEMPR72[14] , 
        \B_DOUT_TEMPR72[13] , \B_DOUT_TEMPR72[12] , 
        \B_DOUT_TEMPR72[11] , \B_DOUT_TEMPR72[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[72][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR2 OR2_64 (.A(\A_DOUT_TEMPR72[31] ), .B(\A_DOUT_TEMPR73[31] ), .Y(
        OR2_64_Y));
    OR4 OR4_558 (.A(\A_DOUT_TEMPR95[0] ), .B(\A_DOUT_TEMPR96[0] ), .C(
        \A_DOUT_TEMPR97[0] ), .D(\A_DOUT_TEMPR98[0] ), .Y(OR4_558_Y));
    OR4 OR4_1904 (.A(\B_DOUT_TEMPR52[39] ), .B(\B_DOUT_TEMPR53[39] ), 
        .C(\B_DOUT_TEMPR54[39] ), .D(\B_DOUT_TEMPR55[39] ), .Y(
        OR4_1904_Y));
    OR4 OR4_2106 (.A(\A_DOUT_TEMPR28[38] ), .B(\A_DOUT_TEMPR29[38] ), 
        .C(\A_DOUT_TEMPR30[38] ), .D(\A_DOUT_TEMPR31[38] ), .Y(
        OR4_2106_Y));
    OR4 OR4_2469 (.A(\A_DOUT_TEMPR68[6] ), .B(\A_DOUT_TEMPR69[6] ), .C(
        \A_DOUT_TEMPR70[6] ), .D(\A_DOUT_TEMPR71[6] ), .Y(OR4_2469_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%50%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R50C2 (
        .A_DOUT({nc6150, nc6151, nc6152, nc6153, nc6154, nc6155, 
        nc6156, nc6157, nc6158, nc6159, nc6160, nc6161, nc6162, nc6163, 
        nc6164, \A_DOUT_TEMPR50[14] , \A_DOUT_TEMPR50[13] , 
        \A_DOUT_TEMPR50[12] , \A_DOUT_TEMPR50[11] , 
        \A_DOUT_TEMPR50[10] }), .B_DOUT({nc6165, nc6166, nc6167, 
        nc6168, nc6169, nc6170, nc6171, nc6172, nc6173, nc6174, nc6175, 
        nc6176, nc6177, nc6178, nc6179, \B_DOUT_TEMPR50[14] , 
        \B_DOUT_TEMPR50[13] , \B_DOUT_TEMPR50[12] , 
        \B_DOUT_TEMPR50[11] , \B_DOUT_TEMPR50[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[50][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2508 (.A(\B_DOUT_TEMPR111[8] ), .B(\B_DOUT_TEMPR112[8] ), 
        .C(\B_DOUT_TEMPR113[8] ), .D(\B_DOUT_TEMPR114[8] ), .Y(
        OR4_2508_Y));
    OR4 OR4_2094 (.A(\B_DOUT_TEMPR32[27] ), .B(\B_DOUT_TEMPR33[27] ), 
        .C(\B_DOUT_TEMPR34[27] ), .D(\B_DOUT_TEMPR35[27] ), .Y(
        OR4_2094_Y));
    OR4 OR4_1748 (.A(OR4_1026_Y), .B(OR4_1912_Y), .C(OR4_1561_Y), .D(
        OR4_34_Y), .Y(OR4_1748_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%31%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R31C4 (
        .A_DOUT({nc6180, nc6181, nc6182, nc6183, nc6184, nc6185, 
        nc6186, nc6187, nc6188, nc6189, nc6190, nc6191, nc6192, nc6193, 
        nc6194, \A_DOUT_TEMPR31[24] , \A_DOUT_TEMPR31[23] , 
        \A_DOUT_TEMPR31[22] , \A_DOUT_TEMPR31[21] , 
        \A_DOUT_TEMPR31[20] }), .B_DOUT({nc6195, nc6196, nc6197, 
        nc6198, nc6199, nc6200, nc6201, nc6202, nc6203, nc6204, nc6205, 
        nc6206, nc6207, nc6208, nc6209, \B_DOUT_TEMPR31[24] , 
        \B_DOUT_TEMPR31[23] , \B_DOUT_TEMPR31[22] , 
        \B_DOUT_TEMPR31[21] , \B_DOUT_TEMPR31[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[31][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_230 (.A(\A_DOUT_TEMPR107[21] ), .B(\A_DOUT_TEMPR108[21] ), 
        .C(\A_DOUT_TEMPR109[21] ), .D(\A_DOUT_TEMPR110[21] ), .Y(
        OR4_230_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%18%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R18C4 (
        .A_DOUT({nc6210, nc6211, nc6212, nc6213, nc6214, nc6215, 
        nc6216, nc6217, nc6218, nc6219, nc6220, nc6221, nc6222, nc6223, 
        nc6224, \A_DOUT_TEMPR18[24] , \A_DOUT_TEMPR18[23] , 
        \A_DOUT_TEMPR18[22] , \A_DOUT_TEMPR18[21] , 
        \A_DOUT_TEMPR18[20] }), .B_DOUT({nc6225, nc6226, nc6227, 
        nc6228, nc6229, nc6230, nc6231, nc6232, nc6233, nc6234, nc6235, 
        nc6236, nc6237, nc6238, nc6239, \B_DOUT_TEMPR18[24] , 
        \B_DOUT_TEMPR18[23] , \B_DOUT_TEMPR18[22] , 
        \B_DOUT_TEMPR18[21] , \B_DOUT_TEMPR18[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[18][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_842 (.A(\B_DOUT_TEMPR24[1] ), .B(\B_DOUT_TEMPR25[1] ), .C(
        \B_DOUT_TEMPR26[1] ), .D(\B_DOUT_TEMPR27[1] ), .Y(OR4_842_Y));
    OR4 OR4_2096 (.A(\B_DOUT_TEMPR40[34] ), .B(\B_DOUT_TEMPR41[34] ), 
        .C(\B_DOUT_TEMPR42[34] ), .D(\B_DOUT_TEMPR43[34] ), .Y(
        OR4_2096_Y));
    OR2 OR2_14 (.A(\B_DOUT_TEMPR72[19] ), .B(\B_DOUT_TEMPR73[19] ), .Y(
        OR2_14_Y));
    OR4 OR4_2432 (.A(\B_DOUT_TEMPR52[30] ), .B(\B_DOUT_TEMPR53[30] ), 
        .C(\B_DOUT_TEMPR54[30] ), .D(\B_DOUT_TEMPR55[30] ), .Y(
        OR4_2432_Y));
    OR4 OR4_1906 (.A(\A_DOUT_TEMPR87[36] ), .B(\A_DOUT_TEMPR88[36] ), 
        .C(\A_DOUT_TEMPR89[36] ), .D(\A_DOUT_TEMPR90[36] ), .Y(
        OR4_1906_Y));
    OR4 OR4_630 (.A(\B_DOUT_TEMPR4[13] ), .B(\B_DOUT_TEMPR5[13] ), .C(
        \B_DOUT_TEMPR6[13] ), .D(\B_DOUT_TEMPR7[13] ), .Y(OR4_630_Y));
    OR4 OR4_2438 (.A(\A_DOUT_TEMPR40[36] ), .B(\A_DOUT_TEMPR41[36] ), 
        .C(\A_DOUT_TEMPR42[36] ), .D(\A_DOUT_TEMPR43[36] ), .Y(
        OR4_2438_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%42%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R42C3 (
        .A_DOUT({nc6240, nc6241, nc6242, nc6243, nc6244, nc6245, 
        nc6246, nc6247, nc6248, nc6249, nc6250, nc6251, nc6252, nc6253, 
        nc6254, \A_DOUT_TEMPR42[19] , \A_DOUT_TEMPR42[18] , 
        \A_DOUT_TEMPR42[17] , \A_DOUT_TEMPR42[16] , 
        \A_DOUT_TEMPR42[15] }), .B_DOUT({nc6255, nc6256, nc6257, 
        nc6258, nc6259, nc6260, nc6261, nc6262, nc6263, nc6264, nc6265, 
        nc6266, nc6267, nc6268, nc6269, \B_DOUT_TEMPR42[19] , 
        \B_DOUT_TEMPR42[18] , \B_DOUT_TEMPR42[17] , 
        \B_DOUT_TEMPR42[16] , \B_DOUT_TEMPR42[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[42][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1432 (.A(\B_DOUT_TEMPR87[33] ), .B(\B_DOUT_TEMPR88[33] ), 
        .C(\B_DOUT_TEMPR89[33] ), .D(\B_DOUT_TEMPR90[33] ), .Y(
        OR4_1432_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%40%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R40C3 (
        .A_DOUT({nc6270, nc6271, nc6272, nc6273, nc6274, nc6275, 
        nc6276, nc6277, nc6278, nc6279, nc6280, nc6281, nc6282, nc6283, 
        nc6284, \A_DOUT_TEMPR40[19] , \A_DOUT_TEMPR40[18] , 
        \A_DOUT_TEMPR40[17] , \A_DOUT_TEMPR40[16] , 
        \A_DOUT_TEMPR40[15] }), .B_DOUT({nc6285, nc6286, nc6287, 
        nc6288, nc6289, nc6290, nc6291, nc6292, nc6293, nc6294, nc6295, 
        nc6296, nc6297, nc6298, nc6299, \B_DOUT_TEMPR40[19] , 
        \B_DOUT_TEMPR40[18] , \B_DOUT_TEMPR40[17] , 
        \B_DOUT_TEMPR40[16] , \B_DOUT_TEMPR40[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[40][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1060 (.A(\A_DOUT_TEMPR32[27] ), .B(\A_DOUT_TEMPR33[27] ), 
        .C(\A_DOUT_TEMPR34[27] ), .D(\A_DOUT_TEMPR35[27] ), .Y(
        OR4_1060_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%118%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R118C1 (
        .A_DOUT({nc6300, nc6301, nc6302, nc6303, nc6304, nc6305, 
        nc6306, nc6307, nc6308, nc6309, nc6310, nc6311, nc6312, nc6313, 
        nc6314, \A_DOUT_TEMPR118[9] , \A_DOUT_TEMPR118[8] , 
        \A_DOUT_TEMPR118[7] , \A_DOUT_TEMPR118[6] , 
        \A_DOUT_TEMPR118[5] }), .B_DOUT({nc6315, nc6316, nc6317, 
        nc6318, nc6319, nc6320, nc6321, nc6322, nc6323, nc6324, nc6325, 
        nc6326, nc6327, nc6328, nc6329, \B_DOUT_TEMPR118[9] , 
        \B_DOUT_TEMPR118[8] , \B_DOUT_TEMPR118[7] , 
        \B_DOUT_TEMPR118[6] , \B_DOUT_TEMPR118[5] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[118][1] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[9], 
        B_DIN[8], B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_3038 (.A(\B_DOUT_TEMPR48[32] ), .B(\B_DOUT_TEMPR49[32] ), 
        .C(\B_DOUT_TEMPR50[32] ), .D(\B_DOUT_TEMPR51[32] ), .Y(
        OR4_3038_Y));
    OR4 OR4_2413 (.A(\A_DOUT_TEMPR52[27] ), .B(\A_DOUT_TEMPR53[27] ), 
        .C(\A_DOUT_TEMPR54[27] ), .D(\A_DOUT_TEMPR55[27] ), .Y(
        OR4_2413_Y));
    OR4 OR4_907 (.A(OR4_1862_Y), .B(OR4_2149_Y), .C(OR4_1790_Y), .D(
        OR4_2162_Y), .Y(OR4_907_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%5%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R5C1 (
        .A_DOUT({nc6330, nc6331, nc6332, nc6333, nc6334, nc6335, 
        nc6336, nc6337, nc6338, nc6339, nc6340, nc6341, nc6342, nc6343, 
        nc6344, \A_DOUT_TEMPR5[9] , \A_DOUT_TEMPR5[8] , 
        \A_DOUT_TEMPR5[7] , \A_DOUT_TEMPR5[6] , \A_DOUT_TEMPR5[5] }), 
        .B_DOUT({nc6345, nc6346, nc6347, nc6348, nc6349, nc6350, 
        nc6351, nc6352, nc6353, nc6354, nc6355, nc6356, nc6357, nc6358, 
        nc6359, \B_DOUT_TEMPR5[9] , \B_DOUT_TEMPR5[8] , 
        \B_DOUT_TEMPR5[7] , \B_DOUT_TEMPR5[6] , \B_DOUT_TEMPR5[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[5][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[1] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[1] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1438 (.A(\B_DOUT_TEMPR75[39] ), .B(\B_DOUT_TEMPR76[39] ), 
        .C(\B_DOUT_TEMPR77[39] ), .D(\B_DOUT_TEMPR78[39] ), .Y(
        OR4_1438_Y));
    OR4 OR4_355 (.A(\B_DOUT_TEMPR111[39] ), .B(\B_DOUT_TEMPR112[39] ), 
        .C(\B_DOUT_TEMPR113[39] ), .D(\B_DOUT_TEMPR114[39] ), .Y(
        OR4_355_Y));
    OR4 OR4_2324 (.A(\A_DOUT_TEMPR28[3] ), .B(\A_DOUT_TEMPR29[3] ), .C(
        \A_DOUT_TEMPR30[3] ), .D(\A_DOUT_TEMPR31[3] ), .Y(OR4_2324_Y));
    OR4 OR4_727 (.A(OR4_286_Y), .B(OR4_95_Y), .C(OR4_994_Y), .D(
        OR4_2147_Y), .Y(OR4_727_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%73%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R73C1 (
        .A_DOUT({nc6360, nc6361, nc6362, nc6363, nc6364, nc6365, 
        nc6366, nc6367, nc6368, nc6369, nc6370, nc6371, nc6372, nc6373, 
        nc6374, \A_DOUT_TEMPR73[9] , \A_DOUT_TEMPR73[8] , 
        \A_DOUT_TEMPR73[7] , \A_DOUT_TEMPR73[6] , \A_DOUT_TEMPR73[5] })
        , .B_DOUT({nc6375, nc6376, nc6377, nc6378, nc6379, nc6380, 
        nc6381, nc6382, nc6383, nc6384, nc6385, nc6386, nc6387, nc6388, 
        nc6389, \B_DOUT_TEMPR73[9] , \B_DOUT_TEMPR73[8] , 
        \B_DOUT_TEMPR73[7] , \B_DOUT_TEMPR73[6] , \B_DOUT_TEMPR73[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[73][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2393 (.A(\B_DOUT_TEMPR79[6] ), .B(\B_DOUT_TEMPR80[6] ), .C(
        \B_DOUT_TEMPR81[6] ), .D(\B_DOUT_TEMPR82[6] ), .Y(OR4_2393_Y));
    OR4 OR4_323 (.A(\A_DOUT_TEMPR60[36] ), .B(\A_DOUT_TEMPR61[36] ), 
        .C(\A_DOUT_TEMPR62[36] ), .D(\A_DOUT_TEMPR63[36] ), .Y(
        OR4_323_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%31%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R31C3 (
        .A_DOUT({nc6390, nc6391, nc6392, nc6393, nc6394, nc6395, 
        nc6396, nc6397, nc6398, nc6399, nc6400, nc6401, nc6402, nc6403, 
        nc6404, \A_DOUT_TEMPR31[19] , \A_DOUT_TEMPR31[18] , 
        \A_DOUT_TEMPR31[17] , \A_DOUT_TEMPR31[16] , 
        \A_DOUT_TEMPR31[15] }), .B_DOUT({nc6405, nc6406, nc6407, 
        nc6408, nc6409, nc6410, nc6411, nc6412, nc6413, nc6414, nc6415, 
        nc6416, nc6417, nc6418, nc6419, \B_DOUT_TEMPR31[19] , 
        \B_DOUT_TEMPR31[18] , \B_DOUT_TEMPR31[17] , 
        \B_DOUT_TEMPR31[16] , \B_DOUT_TEMPR31[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[31][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2360 (.A(\A_DOUT_TEMPR44[34] ), .B(\A_DOUT_TEMPR45[34] ), 
        .C(\A_DOUT_TEMPR46[34] ), .D(\A_DOUT_TEMPR47[34] ), .Y(
        OR4_2360_Y));
    OR4 OR4_2467 (.A(\B_DOUT_TEMPR36[27] ), .B(\B_DOUT_TEMPR37[27] ), 
        .C(\B_DOUT_TEMPR38[27] ), .D(\B_DOUT_TEMPR39[27] ), .Y(
        OR4_2467_Y));
    OR4 OR4_1127 (.A(OR4_1506_Y), .B(OR4_2310_Y), .C(OR2_32_Y), .D(
        \B_DOUT_TEMPR74[26] ), .Y(OR4_1127_Y));
    OR4 OR4_2084 (.A(OR4_960_Y), .B(OR4_395_Y), .C(OR4_1545_Y), .D(
        OR4_1712_Y), .Y(OR4_2084_Y));
    OR4 OR4_728 (.A(\B_DOUT_TEMPR4[39] ), .B(\B_DOUT_TEMPR5[39] ), .C(
        \B_DOUT_TEMPR6[39] ), .D(\B_DOUT_TEMPR7[39] ), .Y(OR4_728_Y));
    OR4 OR4_1624 (.A(\B_DOUT_TEMPR52[37] ), .B(\B_DOUT_TEMPR53[37] ), 
        .C(\B_DOUT_TEMPR54[37] ), .D(\B_DOUT_TEMPR55[37] ), .Y(
        OR4_1624_Y));
    OR4 OR4_2086 (.A(\B_DOUT_TEMPR56[30] ), .B(\B_DOUT_TEMPR57[30] ), 
        .C(\B_DOUT_TEMPR58[30] ), .D(\B_DOUT_TEMPR59[30] ), .Y(
        OR4_2086_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%88%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R88C6 (
        .A_DOUT({nc6420, nc6421, nc6422, nc6423, nc6424, nc6425, 
        nc6426, nc6427, nc6428, nc6429, nc6430, nc6431, nc6432, nc6433, 
        nc6434, \A_DOUT_TEMPR88[34] , \A_DOUT_TEMPR88[33] , 
        \A_DOUT_TEMPR88[32] , \A_DOUT_TEMPR88[31] , 
        \A_DOUT_TEMPR88[30] }), .B_DOUT({nc6435, nc6436, nc6437, 
        nc6438, nc6439, nc6440, nc6441, nc6442, nc6443, nc6444, nc6445, 
        nc6446, nc6447, nc6448, nc6449, \B_DOUT_TEMPR88[34] , 
        \B_DOUT_TEMPR88[33] , \B_DOUT_TEMPR88[32] , 
        \B_DOUT_TEMPR88[31] , \B_DOUT_TEMPR88[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[88][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%118%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R118C3 (
        .A_DOUT({nc6450, nc6451, nc6452, nc6453, nc6454, nc6455, 
        nc6456, nc6457, nc6458, nc6459, nc6460, nc6461, nc6462, nc6463, 
        nc6464, \A_DOUT_TEMPR118[19] , \A_DOUT_TEMPR118[18] , 
        \A_DOUT_TEMPR118[17] , \A_DOUT_TEMPR118[16] , 
        \A_DOUT_TEMPR118[15] }), .B_DOUT({nc6465, nc6466, nc6467, 
        nc6468, nc6469, nc6470, nc6471, nc6472, nc6473, nc6474, nc6475, 
        nc6476, nc6477, nc6478, nc6479, \B_DOUT_TEMPR118[19] , 
        \B_DOUT_TEMPR118[18] , \B_DOUT_TEMPR118[17] , 
        \B_DOUT_TEMPR118[16] , \B_DOUT_TEMPR118[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[118][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_623 (.A(\B_DOUT_TEMPR56[8] ), .B(\B_DOUT_TEMPR57[8] ), .C(
        \B_DOUT_TEMPR58[8] ), .D(\B_DOUT_TEMPR59[8] ), .Y(OR4_623_Y));
    OR4 OR4_2530 (.A(\B_DOUT_TEMPR103[0] ), .B(\B_DOUT_TEMPR104[0] ), 
        .C(\B_DOUT_TEMPR105[0] ), .D(\B_DOUT_TEMPR106[0] ), .Y(
        OR4_2530_Y));
    OR4 OR4_506 (.A(\B_DOUT_TEMPR28[24] ), .B(\B_DOUT_TEMPR29[24] ), 
        .C(\B_DOUT_TEMPR30[24] ), .D(\B_DOUT_TEMPR31[24] ), .Y(
        OR4_506_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%46%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R46C6 (
        .A_DOUT({nc6480, nc6481, nc6482, nc6483, nc6484, nc6485, 
        nc6486, nc6487, nc6488, nc6489, nc6490, nc6491, nc6492, nc6493, 
        nc6494, \A_DOUT_TEMPR46[34] , \A_DOUT_TEMPR46[33] , 
        \A_DOUT_TEMPR46[32] , \A_DOUT_TEMPR46[31] , 
        \A_DOUT_TEMPR46[30] }), .B_DOUT({nc6495, nc6496, nc6497, 
        nc6498, nc6499, nc6500, nc6501, nc6502, nc6503, nc6504, nc6505, 
        nc6506, nc6507, nc6508, nc6509, \B_DOUT_TEMPR46[34] , 
        \B_DOUT_TEMPR46[33] , \B_DOUT_TEMPR46[32] , 
        \B_DOUT_TEMPR46[31] , \B_DOUT_TEMPR46[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[46][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1119 (.A(\A_DOUT_TEMPR56[17] ), .B(\A_DOUT_TEMPR57[17] ), 
        .C(\A_DOUT_TEMPR58[17] ), .D(\A_DOUT_TEMPR59[17] ), .Y(
        OR4_1119_Y));
    OR4 \OR4_A_DOUT[21]  (.A(OR4_225_Y), .B(OR4_2882_Y), .C(OR4_2537_Y)
        , .D(OR4_1474_Y), .Y(A_DOUT[21]));
    OR4 OR4_1530 (.A(\B_DOUT_TEMPR8[2] ), .B(\B_DOUT_TEMPR9[2] ), .C(
        \B_DOUT_TEMPR10[2] ), .D(\B_DOUT_TEMPR11[2] ), .Y(OR4_1530_Y));
    OR4 OR4_98 (.A(OR4_164_Y), .B(OR4_485_Y), .C(OR4_108_Y), .D(
        OR4_505_Y), .Y(OR4_98_Y));
    OR4 OR4_1698 (.A(\B_DOUT_TEMPR91[10] ), .B(\B_DOUT_TEMPR92[10] ), 
        .C(\B_DOUT_TEMPR93[10] ), .D(\B_DOUT_TEMPR94[10] ), .Y(
        OR4_1698_Y));
    OR4 OR4_2383 (.A(\A_DOUT_TEMPR44[3] ), .B(\A_DOUT_TEMPR45[3] ), .C(
        \A_DOUT_TEMPR46[3] ), .D(\A_DOUT_TEMPR47[3] ), .Y(OR4_2383_Y));
    OR4 OR4_1480 (.A(\B_DOUT_TEMPR79[31] ), .B(\B_DOUT_TEMPR80[31] ), 
        .C(\B_DOUT_TEMPR81[31] ), .D(\B_DOUT_TEMPR82[31] ), .Y(
        OR4_1480_Y));
    OR4 OR4_2577 (.A(OR4_2219_Y), .B(OR4_163_Y), .C(OR4_2240_Y), .D(
        OR4_762_Y), .Y(OR4_2577_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%30%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R30C2 (
        .A_DOUT({nc6510, nc6511, nc6512, nc6513, nc6514, nc6515, 
        nc6516, nc6517, nc6518, nc6519, nc6520, nc6521, nc6522, nc6523, 
        nc6524, \A_DOUT_TEMPR30[14] , \A_DOUT_TEMPR30[13] , 
        \A_DOUT_TEMPR30[12] , \A_DOUT_TEMPR30[11] , 
        \A_DOUT_TEMPR30[10] }), .B_DOUT({nc6525, nc6526, nc6527, 
        nc6528, nc6529, nc6530, nc6531, nc6532, nc6533, nc6534, nc6535, 
        nc6536, nc6537, nc6538, nc6539, \B_DOUT_TEMPR30[14] , 
        \B_DOUT_TEMPR30[13] , \B_DOUT_TEMPR30[12] , 
        \B_DOUT_TEMPR30[11] , \B_DOUT_TEMPR30[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[30][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_796 (.A(OR4_1726_Y), .B(OR4_2038_Y), .C(OR4_601_Y), .D(
        OR4_1516_Y), .Y(OR4_796_Y));
    OR4 OR4_850 (.A(\A_DOUT_TEMPR20[12] ), .B(\A_DOUT_TEMPR21[12] ), 
        .C(\A_DOUT_TEMPR22[12] ), .D(\A_DOUT_TEMPR23[12] ), .Y(
        OR4_850_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%14%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R14C7 (
        .A_DOUT({nc6540, nc6541, nc6542, nc6543, nc6544, nc6545, 
        nc6546, nc6547, nc6548, nc6549, nc6550, nc6551, nc6552, nc6553, 
        nc6554, \A_DOUT_TEMPR14[39] , \A_DOUT_TEMPR14[38] , 
        \A_DOUT_TEMPR14[37] , \A_DOUT_TEMPR14[36] , 
        \A_DOUT_TEMPR14[35] }), .B_DOUT({nc6555, nc6556, nc6557, 
        nc6558, nc6559, nc6560, nc6561, nc6562, nc6563, nc6564, nc6565, 
        nc6566, nc6567, nc6568, nc6569, \B_DOUT_TEMPR14[39] , 
        \B_DOUT_TEMPR14[38] , \B_DOUT_TEMPR14[37] , 
        \B_DOUT_TEMPR14[36] , \B_DOUT_TEMPR14[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[14][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1466 (.A(\B_DOUT_TEMPR28[4] ), .B(\B_DOUT_TEMPR29[4] ), .C(
        \B_DOUT_TEMPR30[4] ), .D(\B_DOUT_TEMPR31[4] ), .Y(OR4_1466_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%63%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R63C4 (
        .A_DOUT({nc6570, nc6571, nc6572, nc6573, nc6574, nc6575, 
        nc6576, nc6577, nc6578, nc6579, nc6580, nc6581, nc6582, nc6583, 
        nc6584, \A_DOUT_TEMPR63[24] , \A_DOUT_TEMPR63[23] , 
        \A_DOUT_TEMPR63[22] , \A_DOUT_TEMPR63[21] , 
        \A_DOUT_TEMPR63[20] }), .B_DOUT({nc6585, nc6586, nc6587, 
        nc6588, nc6589, nc6590, nc6591, nc6592, nc6593, nc6594, nc6595, 
        nc6596, nc6597, nc6598, nc6599, \B_DOUT_TEMPR63[24] , 
        \B_DOUT_TEMPR63[23] , \B_DOUT_TEMPR63[22] , 
        \B_DOUT_TEMPR63[21] , \B_DOUT_TEMPR63[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[63][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_550 (.A(\B_DOUT_TEMPR12[35] ), .B(\B_DOUT_TEMPR13[35] ), 
        .C(\B_DOUT_TEMPR14[35] ), .D(\B_DOUT_TEMPR15[35] ), .Y(
        OR4_550_Y));
    OR4 OR4_51 (.A(\B_DOUT_TEMPR87[38] ), .B(\B_DOUT_TEMPR88[38] ), .C(
        \B_DOUT_TEMPR89[38] ), .D(\B_DOUT_TEMPR90[38] ), .Y(OR4_51_Y));
    OR4 OR4_1074 (.A(\A_DOUT_TEMPR103[11] ), .B(\A_DOUT_TEMPR104[11] ), 
        .C(\A_DOUT_TEMPR105[11] ), .D(\A_DOUT_TEMPR106[11] ), .Y(
        OR4_1074_Y));
    OR4 OR4_2159 (.A(OR4_1843_Y), .B(OR4_2142_Y), .C(OR4_1774_Y), .D(
        OR4_2152_Y), .Y(OR4_2159_Y));
    OR4 OR4_1076 (.A(OR4_615_Y), .B(OR4_2104_Y), .C(OR4_2709_Y), .D(
        OR4_2504_Y), .Y(OR4_1076_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%22%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R22C5 (
        .A_DOUT({nc6600, nc6601, nc6602, nc6603, nc6604, nc6605, 
        nc6606, nc6607, nc6608, nc6609, nc6610, nc6611, nc6612, nc6613, 
        nc6614, \A_DOUT_TEMPR22[29] , \A_DOUT_TEMPR22[28] , 
        \A_DOUT_TEMPR22[27] , \A_DOUT_TEMPR22[26] , 
        \A_DOUT_TEMPR22[25] }), .B_DOUT({nc6615, nc6616, nc6617, 
        nc6618, nc6619, nc6620, nc6621, nc6622, nc6623, nc6624, nc6625, 
        nc6626, nc6627, nc6628, nc6629, \B_DOUT_TEMPR22[29] , 
        \B_DOUT_TEMPR22[28] , \B_DOUT_TEMPR22[27] , 
        \B_DOUT_TEMPR22[26] , \B_DOUT_TEMPR22[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[22][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1285 (.A(\B_DOUT_TEMPR79[16] ), .B(\B_DOUT_TEMPR80[16] ), 
        .C(\B_DOUT_TEMPR81[16] ), .D(\B_DOUT_TEMPR82[16] ), .Y(
        OR4_1285_Y));
    OR4 OR4_2504 (.A(\A_DOUT_TEMPR28[30] ), .B(\A_DOUT_TEMPR29[30] ), 
        .C(\A_DOUT_TEMPR30[30] ), .D(\A_DOUT_TEMPR31[30] ), .Y(
        OR4_2504_Y));
    OR4 OR4_1557 (.A(\B_DOUT_TEMPR0[7] ), .B(\B_DOUT_TEMPR1[7] ), .C(
        \B_DOUT_TEMPR2[7] ), .D(\B_DOUT_TEMPR3[7] ), .Y(OR4_1557_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%84%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R84C3 (
        .A_DOUT({nc6630, nc6631, nc6632, nc6633, nc6634, nc6635, 
        nc6636, nc6637, nc6638, nc6639, nc6640, nc6641, nc6642, nc6643, 
        nc6644, \A_DOUT_TEMPR84[19] , \A_DOUT_TEMPR84[18] , 
        \A_DOUT_TEMPR84[17] , \A_DOUT_TEMPR84[16] , 
        \A_DOUT_TEMPR84[15] }), .B_DOUT({nc6645, nc6646, nc6647, 
        nc6648, nc6649, nc6650, nc6651, nc6652, nc6653, nc6654, nc6655, 
        nc6656, nc6657, nc6658, nc6659, \B_DOUT_TEMPR84[19] , 
        \B_DOUT_TEMPR84[18] , \B_DOUT_TEMPR84[17] , 
        \B_DOUT_TEMPR84[16] , \B_DOUT_TEMPR84[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[84][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_754 (.A(OR4_1332_Y), .B(OR4_2764_Y), .C(OR4_2211_Y), .D(
        OR4_625_Y), .Y(OR4_754_Y));
    OR4 OR4_2935 (.A(\A_DOUT_TEMPR24[18] ), .B(\A_DOUT_TEMPR25[18] ), 
        .C(\A_DOUT_TEMPR26[18] ), .D(\A_DOUT_TEMPR27[18] ), .Y(
        OR4_2935_Y));
    OR4 OR4_747 (.A(\B_DOUT_TEMPR24[33] ), .B(\B_DOUT_TEMPR25[33] ), 
        .C(\B_DOUT_TEMPR26[33] ), .D(\B_DOUT_TEMPR27[33] ), .Y(
        OR4_747_Y));
    OR4 OR4_1765 (.A(\B_DOUT_TEMPR91[15] ), .B(\B_DOUT_TEMPR92[15] ), 
        .C(\B_DOUT_TEMPR93[15] ), .D(\B_DOUT_TEMPR94[15] ), .Y(
        OR4_1765_Y));
    OR4 OR4_343 (.A(\A_DOUT_TEMPR68[34] ), .B(\A_DOUT_TEMPR69[34] ), 
        .C(\A_DOUT_TEMPR70[34] ), .D(\A_DOUT_TEMPR71[34] ), .Y(
        OR4_343_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%54%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R54C6 (
        .A_DOUT({nc6660, nc6661, nc6662, nc6663, nc6664, nc6665, 
        nc6666, nc6667, nc6668, nc6669, nc6670, nc6671, nc6672, nc6673, 
        nc6674, \A_DOUT_TEMPR54[34] , \A_DOUT_TEMPR54[33] , 
        \A_DOUT_TEMPR54[32] , \A_DOUT_TEMPR54[31] , 
        \A_DOUT_TEMPR54[30] }), .B_DOUT({nc6675, nc6676, nc6677, 
        nc6678, nc6679, nc6680, nc6681, nc6682, nc6683, nc6684, nc6685, 
        nc6686, nc6687, nc6688, nc6689, \B_DOUT_TEMPR54[34] , 
        \B_DOUT_TEMPR54[33] , \B_DOUT_TEMPR54[32] , 
        \B_DOUT_TEMPR54[31] , \B_DOUT_TEMPR54[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[54][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%22%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R22C1 (
        .A_DOUT({nc6690, nc6691, nc6692, nc6693, nc6694, nc6695, 
        nc6696, nc6697, nc6698, nc6699, nc6700, nc6701, nc6702, nc6703, 
        nc6704, \A_DOUT_TEMPR22[9] , \A_DOUT_TEMPR22[8] , 
        \A_DOUT_TEMPR22[7] , \A_DOUT_TEMPR22[6] , \A_DOUT_TEMPR22[5] })
        , .B_DOUT({nc6705, nc6706, nc6707, nc6708, nc6709, nc6710, 
        nc6711, nc6712, nc6713, nc6714, nc6715, nc6716, nc6717, nc6718, 
        nc6719, \B_DOUT_TEMPR22[9] , \B_DOUT_TEMPR22[8] , 
        \B_DOUT_TEMPR22[7] , \B_DOUT_TEMPR22[6] , \B_DOUT_TEMPR22[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[22][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], 
        A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1935 (.A(OR4_1989_Y), .B(OR4_2829_Y), .C(OR4_1867_Y), .D(
        OR4_1418_Y), .Y(OR4_1935_Y));
    OR4 OR4_591 (.A(\B_DOUT_TEMPR48[6] ), .B(\B_DOUT_TEMPR49[6] ), .C(
        \B_DOUT_TEMPR50[6] ), .D(\B_DOUT_TEMPR51[6] ), .Y(OR4_591_Y));
    OR4 OR4_748 (.A(OR4_1980_Y), .B(OR4_1788_Y), .C(OR4_1728_Y), .D(
        OR4_2230_Y), .Y(OR4_748_Y));
    OR4 OR4_598 (.A(\B_DOUT_TEMPR87[28] ), .B(\B_DOUT_TEMPR88[28] ), 
        .C(\B_DOUT_TEMPR89[28] ), .D(\B_DOUT_TEMPR90[28] ), .Y(
        OR4_598_Y));
    OR4 OR4_2639 (.A(\A_DOUT_TEMPR12[2] ), .B(\A_DOUT_TEMPR13[2] ), .C(
        \A_DOUT_TEMPR14[2] ), .D(\A_DOUT_TEMPR15[2] ), .Y(OR4_2639_Y));
    OR4 OR4_1373 (.A(OR4_101_Y), .B(OR4_1310_Y), .C(OR2_55_Y), .D(
        \B_DOUT_TEMPR74[16] ), .Y(OR4_1373_Y));
    OR4 OR4_2420 (.A(\B_DOUT_TEMPR36[18] ), .B(\B_DOUT_TEMPR37[18] ), 
        .C(\B_DOUT_TEMPR38[18] ), .D(\B_DOUT_TEMPR39[18] ), .Y(
        OR4_2420_Y));
    OR4 OR4_643 (.A(\A_DOUT_TEMPR60[19] ), .B(\A_DOUT_TEMPR61[19] ), 
        .C(\A_DOUT_TEMPR62[19] ), .D(\A_DOUT_TEMPR63[19] ), .Y(
        OR4_643_Y));
    OR4 OR4_1639 (.A(\B_DOUT_TEMPR36[26] ), .B(\B_DOUT_TEMPR37[26] ), 
        .C(\B_DOUT_TEMPR38[26] ), .D(\B_DOUT_TEMPR39[26] ), .Y(
        OR4_1639_Y));
    OR4 OR4_2848 (.A(\A_DOUT_TEMPR48[25] ), .B(\A_DOUT_TEMPR49[25] ), 
        .C(\A_DOUT_TEMPR50[25] ), .D(\A_DOUT_TEMPR51[25] ), .Y(
        OR4_2848_Y));
    OR4 OR4_957 (.A(\A_DOUT_TEMPR44[6] ), .B(\A_DOUT_TEMPR45[6] ), .C(
        \A_DOUT_TEMPR46[6] ), .D(\A_DOUT_TEMPR47[6] ), .Y(OR4_957_Y));
    OR4 OR4_823 (.A(\A_DOUT_TEMPR0[7] ), .B(\A_DOUT_TEMPR1[7] ), .C(
        \A_DOUT_TEMPR2[7] ), .D(\A_DOUT_TEMPR3[7] ), .Y(OR4_823_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%98%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R98C0 (
        .A_DOUT({nc6720, nc6721, nc6722, nc6723, nc6724, nc6725, 
        nc6726, nc6727, nc6728, nc6729, nc6730, nc6731, nc6732, nc6733, 
        nc6734, \A_DOUT_TEMPR98[4] , \A_DOUT_TEMPR98[3] , 
        \A_DOUT_TEMPR98[2] , \A_DOUT_TEMPR98[1] , \A_DOUT_TEMPR98[0] })
        , .B_DOUT({nc6735, nc6736, nc6737, nc6738, nc6739, nc6740, 
        nc6741, nc6742, nc6743, nc6744, nc6745, nc6746, nc6747, nc6748, 
        nc6749, \B_DOUT_TEMPR98[4] , \B_DOUT_TEMPR98[3] , 
        \B_DOUT_TEMPR98[2] , \B_DOUT_TEMPR98[1] , \B_DOUT_TEMPR98[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[98][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2201 (.A(OR4_3015_Y), .B(OR4_1180_Y), .C(OR4_1845_Y), .D(
        OR4_2138_Y), .Y(OR4_2201_Y));
    OR4 OR4_2216 (.A(OR4_1505_Y), .B(OR4_2721_Y), .C(OR2_22_Y), .D(
        \A_DOUT_TEMPR74[19] ), .Y(OR4_2216_Y));
    OR2 OR2_51 (.A(\A_DOUT_TEMPR72[33] ), .B(\A_DOUT_TEMPR73[33] ), .Y(
        OR2_51_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%61%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R61C4 (
        .A_DOUT({nc6750, nc6751, nc6752, nc6753, nc6754, nc6755, 
        nc6756, nc6757, nc6758, nc6759, nc6760, nc6761, nc6762, nc6763, 
        nc6764, \A_DOUT_TEMPR61[24] , \A_DOUT_TEMPR61[23] , 
        \A_DOUT_TEMPR61[22] , \A_DOUT_TEMPR61[21] , 
        \A_DOUT_TEMPR61[20] }), .B_DOUT({nc6765, nc6766, nc6767, 
        nc6768, nc6769, nc6770, nc6771, nc6772, nc6773, nc6774, nc6775, 
        nc6776, nc6777, nc6778, nc6779, \B_DOUT_TEMPR61[24] , 
        \B_DOUT_TEMPR61[23] , \B_DOUT_TEMPR61[22] , 
        \B_DOUT_TEMPR61[21] , \B_DOUT_TEMPR61[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[61][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_689 (.A(OR4_51_Y), .B(OR4_981_Y), .C(OR4_610_Y), .D(
        OR4_2098_Y), .Y(OR4_689_Y));
    OR4 OR4_2278 (.A(\A_DOUT_TEMPR40[6] ), .B(\A_DOUT_TEMPR41[6] ), .C(
        \A_DOUT_TEMPR42[6] ), .D(\A_DOUT_TEMPR43[6] ), .Y(OR4_2278_Y));
    OR4 OR4_2225 (.A(\A_DOUT_TEMPR75[5] ), .B(\A_DOUT_TEMPR76[5] ), .C(
        \A_DOUT_TEMPR77[5] ), .D(\A_DOUT_TEMPR78[5] ), .Y(OR4_2225_Y));
    OR4 OR4_395 (.A(OR4_2186_Y), .B(OR4_2018_Y), .C(OR4_2907_Y), .D(
        OR4_1057_Y), .Y(OR4_395_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%114%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R114C3 (
        .A_DOUT({nc6780, nc6781, nc6782, nc6783, nc6784, nc6785, 
        nc6786, nc6787, nc6788, nc6789, nc6790, nc6791, nc6792, nc6793, 
        nc6794, \A_DOUT_TEMPR114[19] , \A_DOUT_TEMPR114[18] , 
        \A_DOUT_TEMPR114[17] , \A_DOUT_TEMPR114[16] , 
        \A_DOUT_TEMPR114[15] }), .B_DOUT({nc6795, nc6796, nc6797, 
        nc6798, nc6799, nc6800, nc6801, nc6802, nc6803, nc6804, nc6805, 
        nc6806, nc6807, nc6808, nc6809, \B_DOUT_TEMPR114[19] , 
        \B_DOUT_TEMPR114[18] , \B_DOUT_TEMPR114[17] , 
        \B_DOUT_TEMPR114[16] , \B_DOUT_TEMPR114[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[114][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_556 (.A(\A_DOUT_TEMPR83[4] ), .B(\A_DOUT_TEMPR84[4] ), .C(
        \A_DOUT_TEMPR85[4] ), .D(\A_DOUT_TEMPR86[4] ), .Y(OR4_556_Y));
    OR4 OR4_1812 (.A(\B_DOUT_TEMPR4[19] ), .B(\B_DOUT_TEMPR5[19] ), .C(
        \B_DOUT_TEMPR6[19] ), .D(\B_DOUT_TEMPR7[19] ), .Y(OR4_1812_Y));
    OR4 OR4_1620 (.A(\A_DOUT_TEMPR40[25] ), .B(\A_DOUT_TEMPR41[25] ), 
        .C(\A_DOUT_TEMPR42[25] ), .D(\A_DOUT_TEMPR43[25] ), .Y(
        OR4_1620_Y));
    OR4 OR4_170 (.A(\A_DOUT_TEMPR99[11] ), .B(\A_DOUT_TEMPR100[11] ), 
        .C(\A_DOUT_TEMPR101[11] ), .D(\A_DOUT_TEMPR102[11] ), .Y(
        OR4_170_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%71%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R71C2 (
        .A_DOUT({nc6810, nc6811, nc6812, nc6813, nc6814, nc6815, 
        nc6816, nc6817, nc6818, nc6819, nc6820, nc6821, nc6822, nc6823, 
        nc6824, \A_DOUT_TEMPR71[14] , \A_DOUT_TEMPR71[13] , 
        \A_DOUT_TEMPR71[12] , \A_DOUT_TEMPR71[11] , 
        \A_DOUT_TEMPR71[10] }), .B_DOUT({nc6825, nc6826, nc6827, 
        nc6828, nc6829, nc6830, nc6831, nc6832, nc6833, nc6834, nc6835, 
        nc6836, nc6837, nc6838, nc6839, \B_DOUT_TEMPR71[14] , 
        \B_DOUT_TEMPR71[13] , \B_DOUT_TEMPR71[12] , 
        \B_DOUT_TEMPR71[11] , \B_DOUT_TEMPR71[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[71][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1149 (.A(\B_DOUT_TEMPR111[4] ), .B(\B_DOUT_TEMPR112[4] ), 
        .C(\B_DOUT_TEMPR113[4] ), .D(\B_DOUT_TEMPR114[4] ), .Y(
        OR4_1149_Y));
    OR4 OR4_1028 (.A(\B_DOUT_TEMPR79[18] ), .B(\B_DOUT_TEMPR80[18] ), 
        .C(\B_DOUT_TEMPR81[18] ), .D(\B_DOUT_TEMPR82[18] ), .Y(
        OR4_1028_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%104%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R104C1 (
        .A_DOUT({nc6840, nc6841, nc6842, nc6843, nc6844, nc6845, 
        nc6846, nc6847, nc6848, nc6849, nc6850, nc6851, nc6852, nc6853, 
        nc6854, \A_DOUT_TEMPR104[9] , \A_DOUT_TEMPR104[8] , 
        \A_DOUT_TEMPR104[7] , \A_DOUT_TEMPR104[6] , 
        \A_DOUT_TEMPR104[5] }), .B_DOUT({nc6855, nc6856, nc6857, 
        nc6858, nc6859, nc6860, nc6861, nc6862, nc6863, nc6864, nc6865, 
        nc6866, nc6867, nc6868, nc6869, \B_DOUT_TEMPR104[9] , 
        \B_DOUT_TEMPR104[8] , \B_DOUT_TEMPR104[7] , 
        \B_DOUT_TEMPR104[6] , \B_DOUT_TEMPR104[5] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[104][1] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[9], 
        B_DIN[8], B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_983 (.A(OR4_260_Y), .B(OR4_2637_Y), .C(OR2_37_Y), .D(
        \B_DOUT_TEMPR74[6] ), .Y(OR4_983_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%61%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R61C3 (
        .A_DOUT({nc6870, nc6871, nc6872, nc6873, nc6874, nc6875, 
        nc6876, nc6877, nc6878, nc6879, nc6880, nc6881, nc6882, nc6883, 
        nc6884, \A_DOUT_TEMPR61[19] , \A_DOUT_TEMPR61[18] , 
        \A_DOUT_TEMPR61[17] , \A_DOUT_TEMPR61[16] , 
        \A_DOUT_TEMPR61[15] }), .B_DOUT({nc6885, nc6886, nc6887, 
        nc6888, nc6889, nc6890, nc6891, nc6892, nc6893, nc6894, nc6895, 
        nc6896, nc6897, nc6898, nc6899, \B_DOUT_TEMPR61[19] , 
        \B_DOUT_TEMPR61[18] , \B_DOUT_TEMPR61[17] , 
        \B_DOUT_TEMPR61[16] , \B_DOUT_TEMPR61[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[61][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_612 (.A(OR4_2458_Y), .B(OR4_2742_Y), .C(OR4_367_Y), .D(
        OR4_671_Y), .Y(OR4_612_Y));
    OR4 OR4_122 (.A(\B_DOUT_TEMPR12[36] ), .B(\B_DOUT_TEMPR13[36] ), 
        .C(\B_DOUT_TEMPR14[36] ), .D(\B_DOUT_TEMPR15[36] ), .Y(
        OR4_122_Y));
    OR4 OR4_1258 (.A(\A_DOUT_TEMPR68[7] ), .B(\A_DOUT_TEMPR69[7] ), .C(
        \A_DOUT_TEMPR70[7] ), .D(\A_DOUT_TEMPR71[7] ), .Y(OR4_1258_Y));
    OR4 OR4_678 (.A(\B_DOUT_TEMPR87[9] ), .B(\B_DOUT_TEMPR88[9] ), .C(
        \B_DOUT_TEMPR89[9] ), .D(\B_DOUT_TEMPR90[9] ), .Y(OR4_678_Y));
    OR4 OR4_2064 (.A(OR4_2510_Y), .B(OR4_1184_Y), .C(OR4_1791_Y), .D(
        OR4_1009_Y), .Y(OR4_2064_Y));
    OR4 OR4_1899 (.A(\B_DOUT_TEMPR4[8] ), .B(\B_DOUT_TEMPR5[8] ), .C(
        \B_DOUT_TEMPR6[8] ), .D(\B_DOUT_TEMPR7[8] ), .Y(OR4_1899_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%34%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R34C6 (
        .A_DOUT({nc6900, nc6901, nc6902, nc6903, nc6904, nc6905, 
        nc6906, nc6907, nc6908, nc6909, nc6910, nc6911, nc6912, nc6913, 
        nc6914, \A_DOUT_TEMPR34[34] , \A_DOUT_TEMPR34[33] , 
        \A_DOUT_TEMPR34[32] , \A_DOUT_TEMPR34[31] , 
        \A_DOUT_TEMPR34[30] }), .B_DOUT({nc6915, nc6916, nc6917, 
        nc6918, nc6919, nc6920, nc6921, nc6922, nc6923, nc6924, nc6925, 
        nc6926, nc6927, nc6928, nc6929, \B_DOUT_TEMPR34[34] , 
        \B_DOUT_TEMPR34[33] , \B_DOUT_TEMPR34[32] , 
        \B_DOUT_TEMPR34[31] , \B_DOUT_TEMPR34[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[34][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1686 (.A(\A_DOUT_TEMPR83[23] ), .B(\A_DOUT_TEMPR84[23] ), 
        .C(\A_DOUT_TEMPR85[23] ), .D(\A_DOUT_TEMPR86[23] ), .Y(
        OR4_1686_Y));
    OR4 OR4_2066 (.A(\B_DOUT_TEMPR0[14] ), .B(\B_DOUT_TEMPR1[14] ), .C(
        \B_DOUT_TEMPR2[14] ), .D(\B_DOUT_TEMPR3[14] ), .Y(OR4_2066_Y));
    OR4 OR4_1180 (.A(\B_DOUT_TEMPR36[37] ), .B(\B_DOUT_TEMPR37[37] ), 
        .C(\B_DOUT_TEMPR38[37] ), .D(\B_DOUT_TEMPR39[37] ), .Y(
        OR4_1180_Y));
    OR4 OR4_925 (.A(OR4_2811_Y), .B(OR4_1986_Y), .C(OR4_1422_Y), .D(
        OR4_896_Y), .Y(OR4_925_Y));
    OR4 OR4_1613 (.A(\A_DOUT_TEMPR115[6] ), .B(\A_DOUT_TEMPR116[6] ), 
        .C(\A_DOUT_TEMPR117[6] ), .D(\A_DOUT_TEMPR118[6] ), .Y(
        OR4_1613_Y));
    OR4 OR4_425 (.A(\A_DOUT_TEMPR12[36] ), .B(\A_DOUT_TEMPR13[36] ), 
        .C(\A_DOUT_TEMPR14[36] ), .D(\A_DOUT_TEMPR15[36] ), .Y(
        OR4_425_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%118%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R118C6 (
        .A_DOUT({nc6930, nc6931, nc6932, nc6933, nc6934, nc6935, 
        nc6936, nc6937, nc6938, nc6939, nc6940, nc6941, nc6942, nc6943, 
        nc6944, \A_DOUT_TEMPR118[34] , \A_DOUT_TEMPR118[33] , 
        \A_DOUT_TEMPR118[32] , \A_DOUT_TEMPR118[31] , 
        \A_DOUT_TEMPR118[30] }), .B_DOUT({nc6945, nc6946, nc6947, 
        nc6948, nc6949, nc6950, nc6951, nc6952, nc6953, nc6954, nc6955, 
        nc6956, nc6957, nc6958, nc6959, \B_DOUT_TEMPR118[34] , 
        \B_DOUT_TEMPR118[33] , \B_DOUT_TEMPR118[32] , 
        \B_DOUT_TEMPR118[31] , \B_DOUT_TEMPR118[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[118][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2852 (.A(OR4_307_Y), .B(OR4_1509_Y), .C(OR2_65_Y), .D(
        \A_DOUT_TEMPR74[11] ), .Y(OR4_2852_Y));
    OR4 OR4_890 (.A(\B_DOUT_TEMPR60[5] ), .B(\B_DOUT_TEMPR61[5] ), .C(
        \B_DOUT_TEMPR62[5] ), .D(\B_DOUT_TEMPR63[5] ), .Y(OR4_890_Y));
    OR4 OR4_2748 (.A(\B_DOUT_TEMPR24[24] ), .B(\B_DOUT_TEMPR25[24] ), 
        .C(\B_DOUT_TEMPR26[24] ), .D(\B_DOUT_TEMPR27[24] ), .Y(
        OR4_2748_Y));
    OR4 OR4_2816 (.A(\B_DOUT_TEMPR4[28] ), .B(\B_DOUT_TEMPR5[28] ), .C(
        \B_DOUT_TEMPR6[28] ), .D(\B_DOUT_TEMPR7[28] ), .Y(OR4_2816_Y));
    OR4 OR4_1919 (.A(OR4_2118_Y), .B(OR4_741_Y), .C(OR4_119_Y), .D(
        OR4_2492_Y), .Y(OR4_1919_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%95%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R95C0 (
        .A_DOUT({nc6960, nc6961, nc6962, nc6963, nc6964, nc6965, 
        nc6966, nc6967, nc6968, nc6969, nc6970, nc6971, nc6972, nc6973, 
        nc6974, \A_DOUT_TEMPR95[4] , \A_DOUT_TEMPR95[3] , 
        \A_DOUT_TEMPR95[2] , \A_DOUT_TEMPR95[1] , \A_DOUT_TEMPR95[0] })
        , .B_DOUT({nc6975, nc6976, nc6977, nc6978, nc6979, nc6980, 
        nc6981, nc6982, nc6983, nc6984, nc6985, nc6986, nc6987, nc6988, 
        nc6989, \B_DOUT_TEMPR95[4] , \B_DOUT_TEMPR95[3] , 
        \B_DOUT_TEMPR95[2] , \B_DOUT_TEMPR95[1] , \B_DOUT_TEMPR95[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[95][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_78 (.A(\B_DOUT_TEMPR4[17] ), .B(\B_DOUT_TEMPR5[17] ), .C(
        \B_DOUT_TEMPR6[17] ), .D(\B_DOUT_TEMPR7[17] ), .Y(OR4_78_Y));
    OR4 OR4_590 (.A(\A_DOUT_TEMPR12[6] ), .B(\A_DOUT_TEMPR13[6] ), .C(
        \A_DOUT_TEMPR14[6] ), .D(\A_DOUT_TEMPR15[6] ), .Y(OR4_590_Y));
    OR4 OR4_971 (.A(\B_DOUT_TEMPR91[6] ), .B(\B_DOUT_TEMPR92[6] ), .C(
        \B_DOUT_TEMPR93[6] ), .D(\B_DOUT_TEMPR94[6] ), .Y(OR4_971_Y));
    OR4 OR4_1191 (.A(\A_DOUT_TEMPR111[19] ), .B(\A_DOUT_TEMPR112[19] ), 
        .C(\A_DOUT_TEMPR113[19] ), .D(\A_DOUT_TEMPR114[19] ), .Y(
        OR4_1191_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%60%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R60C2 (
        .A_DOUT({nc6990, nc6991, nc6992, nc6993, nc6994, nc6995, 
        nc6996, nc6997, nc6998, nc6999, nc7000, nc7001, nc7002, nc7003, 
        nc7004, \A_DOUT_TEMPR60[14] , \A_DOUT_TEMPR60[13] , 
        \A_DOUT_TEMPR60[12] , \A_DOUT_TEMPR60[11] , 
        \A_DOUT_TEMPR60[10] }), .B_DOUT({nc7005, nc7006, nc7007, 
        nc7008, nc7009, nc7010, nc7011, nc7012, nc7013, nc7014, nc7015, 
        nc7016, nc7017, nc7018, nc7019, \B_DOUT_TEMPR60[14] , 
        \B_DOUT_TEMPR60[13] , \B_DOUT_TEMPR60[12] , 
        \B_DOUT_TEMPR60[11] , \B_DOUT_TEMPR60[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[60][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_843 (.A(\A_DOUT_TEMPR36[28] ), .B(\A_DOUT_TEMPR37[28] ), 
        .C(\A_DOUT_TEMPR38[28] ), .D(\A_DOUT_TEMPR39[28] ), .Y(
        OR4_843_Y));
    OR4 OR4_2363 (.A(\A_DOUT_TEMPR60[5] ), .B(\A_DOUT_TEMPR61[5] ), .C(
        \A_DOUT_TEMPR62[5] ), .D(\A_DOUT_TEMPR63[5] ), .Y(OR4_2363_Y));
    OR4 OR4_1566 (.A(\B_DOUT_TEMPR52[5] ), .B(\B_DOUT_TEMPR53[5] ), .C(
        \B_DOUT_TEMPR54[5] ), .D(\B_DOUT_TEMPR55[5] ), .Y(OR4_1566_Y));
    OR4 OR4_100 (.A(\A_DOUT_TEMPR60[25] ), .B(\A_DOUT_TEMPR61[25] ), 
        .C(\A_DOUT_TEMPR62[25] ), .D(\A_DOUT_TEMPR63[25] ), .Y(
        OR4_100_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%13%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R13C4 (
        .A_DOUT({nc7020, nc7021, nc7022, nc7023, nc7024, nc7025, 
        nc7026, nc7027, nc7028, nc7029, nc7030, nc7031, nc7032, nc7033, 
        nc7034, \A_DOUT_TEMPR13[24] , \A_DOUT_TEMPR13[23] , 
        \A_DOUT_TEMPR13[22] , \A_DOUT_TEMPR13[21] , 
        \A_DOUT_TEMPR13[20] }), .B_DOUT({nc7035, nc7036, nc7037, 
        nc7038, nc7039, nc7040, nc7041, nc7042, nc7043, nc7044, nc7045, 
        nc7046, nc7047, nc7048, nc7049, \B_DOUT_TEMPR13[24] , 
        \B_DOUT_TEMPR13[23] , \B_DOUT_TEMPR13[22] , 
        \B_DOUT_TEMPR13[21] , \B_DOUT_TEMPR13[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[13][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2037 (.A(OR4_2976_Y), .B(OR4_2800_Y), .C(OR4_2745_Y), .D(
        OR4_2715_Y), .Y(OR4_2037_Y));
    OR4 OR4_1095 (.A(OR4_1537_Y), .B(OR4_1837_Y), .C(OR4_1467_Y), .D(
        OR4_1860_Y), .Y(OR4_1095_Y));
    OR4 OR4_1124 (.A(\B_DOUT_TEMPR8[34] ), .B(\B_DOUT_TEMPR9[34] ), .C(
        \B_DOUT_TEMPR10[34] ), .D(\B_DOUT_TEMPR11[34] ), .Y(OR4_1124_Y)
        );
    OR4 \OR4_A_DOUT[38]  (.A(OR4_1158_Y), .B(OR4_421_Y), .C(OR4_2909_Y)
        , .D(OR4_265_Y), .Y(A_DOUT[38]));
    OR4 OR4_794 (.A(\A_DOUT_TEMPR0[38] ), .B(\A_DOUT_TEMPR1[38] ), .C(
        \A_DOUT_TEMPR2[38] ), .D(\A_DOUT_TEMPR3[38] ), .Y(OR4_794_Y));
    OR4 OR4_2339 (.A(\A_DOUT_TEMPR75[36] ), .B(\A_DOUT_TEMPR76[36] ), 
        .C(\A_DOUT_TEMPR77[36] ), .D(\A_DOUT_TEMPR78[36] ), .Y(
        OR4_2339_Y));
    OR4 OR4_1767 (.A(\A_DOUT_TEMPR107[18] ), .B(\A_DOUT_TEMPR108[18] ), 
        .C(\A_DOUT_TEMPR109[18] ), .D(\A_DOUT_TEMPR110[18] ), .Y(
        OR4_1767_Y));
    OR4 OR4_3017 (.A(\B_DOUT_TEMPR91[34] ), .B(\B_DOUT_TEMPR92[34] ), 
        .C(\B_DOUT_TEMPR93[34] ), .D(\B_DOUT_TEMPR94[34] ), .Y(
        OR4_3017_Y));
    OR4 OR4_56 (.A(\A_DOUT_TEMPR52[8] ), .B(\A_DOUT_TEMPR53[8] ), .C(
        \A_DOUT_TEMPR54[8] ), .D(\A_DOUT_TEMPR55[8] ), .Y(OR4_56_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%46%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R46C0 (
        .A_DOUT({nc7050, nc7051, nc7052, nc7053, nc7054, nc7055, 
        nc7056, nc7057, nc7058, nc7059, nc7060, nc7061, nc7062, nc7063, 
        nc7064, \A_DOUT_TEMPR46[4] , \A_DOUT_TEMPR46[3] , 
        \A_DOUT_TEMPR46[2] , \A_DOUT_TEMPR46[1] , \A_DOUT_TEMPR46[0] })
        , .B_DOUT({nc7065, nc7066, nc7067, nc7068, nc7069, nc7070, 
        nc7071, nc7072, nc7073, nc7074, nc7075, nc7076, nc7077, nc7078, 
        nc7079, \B_DOUT_TEMPR46[4] , \B_DOUT_TEMPR46[3] , 
        \B_DOUT_TEMPR46[2] , \B_DOUT_TEMPR46[1] , \B_DOUT_TEMPR46[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[46][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2237 (.A(\B_DOUT_TEMPR56[6] ), .B(\B_DOUT_TEMPR57[6] ), .C(
        \B_DOUT_TEMPR58[6] ), .D(\B_DOUT_TEMPR59[6] ), .Y(OR4_2237_Y));
    OR4 OR4_1561 (.A(\B_DOUT_TEMPR95[39] ), .B(\B_DOUT_TEMPR96[39] ), 
        .C(\B_DOUT_TEMPR97[39] ), .D(\B_DOUT_TEMPR98[39] ), .Y(
        OR4_1561_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%72%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R72C3 (
        .A_DOUT({nc7080, nc7081, nc7082, nc7083, nc7084, nc7085, 
        nc7086, nc7087, nc7088, nc7089, nc7090, nc7091, nc7092, nc7093, 
        nc7094, \A_DOUT_TEMPR72[19] , \A_DOUT_TEMPR72[18] , 
        \A_DOUT_TEMPR72[17] , \A_DOUT_TEMPR72[16] , 
        \A_DOUT_TEMPR72[15] }), .B_DOUT({nc7095, nc7096, nc7097, 
        nc7098, nc7099, nc7100, nc7101, nc7102, nc7103, nc7104, nc7105, 
        nc7106, nc7107, nc7108, nc7109, \B_DOUT_TEMPR72[19] , 
        \B_DOUT_TEMPR72[18] , \B_DOUT_TEMPR72[17] , 
        \B_DOUT_TEMPR72[16] , \B_DOUT_TEMPR72[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[72][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1037 (.A(\A_DOUT_TEMPR0[9] ), .B(\A_DOUT_TEMPR1[9] ), .C(
        \A_DOUT_TEMPR2[9] ), .D(\A_DOUT_TEMPR3[9] ), .Y(OR4_1037_Y));
    OR4 OR4_1339 (.A(\A_DOUT_TEMPR28[4] ), .B(\A_DOUT_TEMPR29[4] ), .C(
        \A_DOUT_TEMPR30[4] ), .D(\A_DOUT_TEMPR31[4] ), .Y(OR4_1339_Y));
    OR4 OR4_1714 (.A(\B_DOUT_TEMPR64[3] ), .B(\B_DOUT_TEMPR65[3] ), .C(
        \B_DOUT_TEMPR66[3] ), .D(\B_DOUT_TEMPR67[3] ), .Y(OR4_1714_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%70%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R70C3 (
        .A_DOUT({nc7110, nc7111, nc7112, nc7113, nc7114, nc7115, 
        nc7116, nc7117, nc7118, nc7119, nc7120, nc7121, nc7122, nc7123, 
        nc7124, \A_DOUT_TEMPR70[19] , \A_DOUT_TEMPR70[18] , 
        \A_DOUT_TEMPR70[17] , \A_DOUT_TEMPR70[16] , 
        \A_DOUT_TEMPR70[15] }), .B_DOUT({nc7125, nc7126, nc7127, 
        nc7128, nc7129, nc7130, nc7131, nc7132, nc7133, nc7134, nc7135, 
        nc7136, nc7137, nc7138, nc7139, \B_DOUT_TEMPR70[19] , 
        \B_DOUT_TEMPR70[18] , \B_DOUT_TEMPR70[17] , 
        \B_DOUT_TEMPR70[16] , \B_DOUT_TEMPR70[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[70][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2653 (.A(\A_DOUT_TEMPR111[15] ), .B(\A_DOUT_TEMPR112[15] ), 
        .C(\A_DOUT_TEMPR113[15] ), .D(\A_DOUT_TEMPR114[15] ), .Y(
        OR4_2653_Y));
    OR4 OR4_1237 (.A(OR4_2062_Y), .B(OR4_2557_Y), .C(OR4_206_Y), .D(
        OR4_514_Y), .Y(OR4_1237_Y));
    OR4 OR4_2959 (.A(OR4_2841_Y), .B(OR4_614_Y), .C(OR4_276_Y), .D(
        OR4_2045_Y), .Y(OR4_2959_Y));
    OR4 OR4_2626 (.A(\B_DOUT_TEMPR36[7] ), .B(\B_DOUT_TEMPR37[7] ), .C(
        \B_DOUT_TEMPR38[7] ), .D(\B_DOUT_TEMPR39[7] ), .Y(OR4_2626_Y));
    OR4 OR4_1411 (.A(OR4_407_Y), .B(OR4_422_Y), .C(OR4_1140_Y), .D(
        OR4_1420_Y), .Y(OR4_1411_Y));
    OR4 OR4_2930 (.A(\A_DOUT_TEMPR28[12] ), .B(\A_DOUT_TEMPR29[12] ), 
        .C(\A_DOUT_TEMPR30[12] ), .D(\A_DOUT_TEMPR31[12] ), .Y(
        OR4_2930_Y));
    OR4 \OR4_B_DOUT[0]  (.A(OR4_511_Y), .B(OR4_1909_Y), .C(OR4_2975_Y), 
        .D(OR4_2808_Y), .Y(B_DOUT[0]));
    OR4 OR4_608 (.A(\B_DOUT_TEMPR44[0] ), .B(\B_DOUT_TEMPR45[0] ), .C(
        \B_DOUT_TEMPR46[0] ), .D(\B_DOUT_TEMPR47[0] ), .Y(OR4_608_Y));
    OR4 OR4_2120 (.A(OR4_1346_Y), .B(OR4_658_Y), .C(OR4_2584_Y), .D(
        OR4_679_Y), .Y(OR4_2120_Y));
    OR4 OR4_2710 (.A(\B_DOUT_TEMPR60[7] ), .B(\B_DOUT_TEMPR61[7] ), .C(
        \B_DOUT_TEMPR62[7] ), .D(\B_DOUT_TEMPR63[7] ), .Y(OR4_2710_Y));
    OR4 OR4_1897 (.A(\A_DOUT_TEMPR32[8] ), .B(\A_DOUT_TEMPR33[8] ), .C(
        \A_DOUT_TEMPR34[8] ), .D(\A_DOUT_TEMPR35[8] ), .Y(OR4_1897_Y));
    OR4 OR4_142 (.A(\A_DOUT_TEMPR79[20] ), .B(\A_DOUT_TEMPR80[20] ), 
        .C(\A_DOUT_TEMPR81[20] ), .D(\A_DOUT_TEMPR82[20] ), .Y(
        OR4_142_Y));
    OR4 OR4_1930 (.A(\A_DOUT_TEMPR32[21] ), .B(\A_DOUT_TEMPR33[21] ), 
        .C(\A_DOUT_TEMPR34[21] ), .D(\A_DOUT_TEMPR35[21] ), .Y(
        OR4_1930_Y));
    OR4 OR4_997 (.A(\B_DOUT_TEMPR115[26] ), .B(\B_DOUT_TEMPR116[26] ), 
        .C(\B_DOUT_TEMPR117[26] ), .D(\B_DOUT_TEMPR118[26] ), .Y(
        OR4_997_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%76%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R76C6 (
        .A_DOUT({nc7140, nc7141, nc7142, nc7143, nc7144, nc7145, 
        nc7146, nc7147, nc7148, nc7149, nc7150, nc7151, nc7152, nc7153, 
        nc7154, \A_DOUT_TEMPR76[34] , \A_DOUT_TEMPR76[33] , 
        \A_DOUT_TEMPR76[32] , \A_DOUT_TEMPR76[31] , 
        \A_DOUT_TEMPR76[30] }), .B_DOUT({nc7155, nc7156, nc7157, 
        nc7158, nc7159, nc7160, nc7161, nc7162, nc7163, nc7164, nc7165, 
        nc7166, nc7167, nc7168, nc7169, \B_DOUT_TEMPR76[34] , 
        \B_DOUT_TEMPR76[33] , \B_DOUT_TEMPR76[32] , 
        \B_DOUT_TEMPR76[31] , \B_DOUT_TEMPR76[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[76][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1825 (.A(OR4_680_Y), .B(OR4_135_Y), .C(OR4_1312_Y), .D(
        OR4_1468_Y), .Y(OR4_1825_Y));
    OR4 OR4_974 (.A(OR4_454_Y), .B(OR4_1236_Y), .C(OR4_776_Y), .D(
        OR4_2452_Y), .Y(OR4_974_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%82%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R82C6 (
        .A_DOUT({nc7170, nc7171, nc7172, nc7173, nc7174, nc7175, 
        nc7176, nc7177, nc7178, nc7179, nc7180, nc7181, nc7182, nc7183, 
        nc7184, \A_DOUT_TEMPR82[34] , \A_DOUT_TEMPR82[33] , 
        \A_DOUT_TEMPR82[32] , \A_DOUT_TEMPR82[31] , 
        \A_DOUT_TEMPR82[30] }), .B_DOUT({nc7185, nc7186, nc7187, 
        nc7188, nc7189, nc7190, nc7191, nc7192, nc7193, nc7194, nc7195, 
        nc7196, nc7197, nc7198, nc7199, \B_DOUT_TEMPR82[34] , 
        \B_DOUT_TEMPR82[33] , \B_DOUT_TEMPR82[32] , 
        \B_DOUT_TEMPR82[31] , \B_DOUT_TEMPR82[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[82][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2198 (.A(OR4_964_Y), .B(OR4_2937_Y), .C(OR4_1530_Y), .D(
        OR4_2521_Y), .Y(OR4_2198_Y));
    OR4 OR4_1842 (.A(OR4_1045_Y), .B(OR4_50_Y), .C(OR4_241_Y), .D(
        OR4_59_Y), .Y(OR4_1842_Y));
    OR4 OR4_901 (.A(OR4_1108_Y), .B(OR4_1632_Y), .C(OR4_2260_Y), .D(
        OR4_1456_Y), .Y(OR4_901_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%99%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R99C1 (
        .A_DOUT({nc7200, nc7201, nc7202, nc7203, nc7204, nc7205, 
        nc7206, nc7207, nc7208, nc7209, nc7210, nc7211, nc7212, nc7213, 
        nc7214, \A_DOUT_TEMPR99[9] , \A_DOUT_TEMPR99[8] , 
        \A_DOUT_TEMPR99[7] , \A_DOUT_TEMPR99[6] , \A_DOUT_TEMPR99[5] })
        , .B_DOUT({nc7215, nc7216, nc7217, nc7218, nc7219, nc7220, 
        nc7221, nc7222, nc7223, nc7224, nc7225, nc7226, nc7227, nc7228, 
        nc7229, \B_DOUT_TEMPR99[9] , \B_DOUT_TEMPR99[8] , 
        \B_DOUT_TEMPR99[7] , \B_DOUT_TEMPR99[6] , \B_DOUT_TEMPR99[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[99][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_945 (.A(OR4_2525_Y), .B(OR4_382_Y), .C(OR4_1152_Y), .D(
        OR4_2677_Y), .Y(OR4_945_Y));
    OR4 OR4_445 (.A(\A_DOUT_TEMPR95[32] ), .B(\A_DOUT_TEMPR96[32] ), 
        .C(\A_DOUT_TEMPR97[32] ), .D(\A_DOUT_TEMPR98[32] ), .Y(
        OR4_445_Y));
    OR4 OR4_2754 (.A(OR4_175_Y), .B(OR4_268_Y), .C(OR4_1747_Y), .D(
        OR4_270_Y), .Y(OR4_2754_Y));
    OR4 OR4_2732 (.A(\B_DOUT_TEMPR32[28] ), .B(\B_DOUT_TEMPR33[28] ), 
        .C(\B_DOUT_TEMPR34[28] ), .D(\B_DOUT_TEMPR35[28] ), .Y(
        OR4_2732_Y));
    OR4 \OR4_A_DOUT[15]  (.A(OR4_2901_Y), .B(OR4_2767_Y), .C(
        OR4_1913_Y), .D(OR4_2536_Y), .Y(A_DOUT[15]));
    OR4 OR4_596 (.A(\A_DOUT_TEMPR56[21] ), .B(\A_DOUT_TEMPR57[21] ), 
        .C(\A_DOUT_TEMPR58[21] ), .D(\A_DOUT_TEMPR59[21] ), .Y(
        OR4_596_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%89%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R89C0 (
        .A_DOUT({nc7230, nc7231, nc7232, nc7233, nc7234, nc7235, 
        nc7236, nc7237, nc7238, nc7239, nc7240, nc7241, nc7242, nc7243, 
        nc7244, \A_DOUT_TEMPR89[4] , \A_DOUT_TEMPR89[3] , 
        \A_DOUT_TEMPR89[2] , \A_DOUT_TEMPR89[1] , \A_DOUT_TEMPR89[0] })
        , .B_DOUT({nc7245, nc7246, nc7247, nc7248, nc7249, nc7250, 
        nc7251, nc7252, nc7253, nc7254, nc7255, nc7256, nc7257, nc7258, 
        nc7259, \B_DOUT_TEMPR89[4] , \B_DOUT_TEMPR89[3] , 
        \B_DOUT_TEMPR89[2] , \B_DOUT_TEMPR89[1] , \B_DOUT_TEMPR89[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[89][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%11%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R11C4 (
        .A_DOUT({nc7260, nc7261, nc7262, nc7263, nc7264, nc7265, 
        nc7266, nc7267, nc7268, nc7269, nc7270, nc7271, nc7272, nc7273, 
        nc7274, \A_DOUT_TEMPR11[24] , \A_DOUT_TEMPR11[23] , 
        \A_DOUT_TEMPR11[22] , \A_DOUT_TEMPR11[21] , 
        \A_DOUT_TEMPR11[20] }), .B_DOUT({nc7275, nc7276, nc7277, 
        nc7278, nc7279, nc7280, nc7281, nc7282, nc7283, nc7284, nc7285, 
        nc7286, nc7287, nc7288, nc7289, \B_DOUT_TEMPR11[24] , 
        \B_DOUT_TEMPR11[23] , \B_DOUT_TEMPR11[22] , 
        \B_DOUT_TEMPR11[21] , \B_DOUT_TEMPR11[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[11][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2451 (.A(OR4_3007_Y), .B(OR4_2161_Y), .C(OR4_1176_Y), .D(
        OR4_1450_Y), .Y(OR4_2451_Y));
    OR2 OR2_56 (.A(\B_DOUT_TEMPR72[18] ), .B(\B_DOUT_TEMPR73[18] ), .Y(
        OR2_56_Y));
    OR4 OR4_1732 (.A(OR4_563_Y), .B(OR4_2780_Y), .C(OR4_1209_Y), .D(
        OR4_2782_Y), .Y(OR4_1732_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENB[0]  (.A(B_WBYTE_EN[0]), .B(
        B_WEN), .Y(\WBYTEENB[0] ));
    OR4 OR4_1914 (.A(\A_DOUT_TEMPR12[17] ), .B(\A_DOUT_TEMPR13[17] ), 
        .C(\A_DOUT_TEMPR14[17] ), .D(\A_DOUT_TEMPR15[17] ), .Y(
        OR4_1914_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%99%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R99C2 (
        .A_DOUT({nc7290, nc7291, nc7292, nc7293, nc7294, nc7295, 
        nc7296, nc7297, nc7298, nc7299, nc7300, nc7301, nc7302, nc7303, 
        nc7304, \A_DOUT_TEMPR99[14] , \A_DOUT_TEMPR99[13] , 
        \A_DOUT_TEMPR99[12] , \A_DOUT_TEMPR99[11] , 
        \A_DOUT_TEMPR99[10] }), .B_DOUT({nc7305, nc7306, nc7307, 
        nc7308, nc7309, nc7310, nc7311, nc7312, nc7313, nc7314, nc7315, 
        nc7316, nc7317, nc7318, nc7319, \B_DOUT_TEMPR99[14] , 
        \B_DOUT_TEMPR99[13] , \B_DOUT_TEMPR99[12] , 
        \B_DOUT_TEMPR99[11] , \B_DOUT_TEMPR99[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[99][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1983 (.A(OR4_1325_Y), .B(OR4_473_Y), .C(OR4_1953_Y), .D(
        OR4_475_Y), .Y(OR4_1983_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%95%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R95C1 (
        .A_DOUT({nc7320, nc7321, nc7322, nc7323, nc7324, nc7325, 
        nc7326, nc7327, nc7328, nc7329, nc7330, nc7331, nc7332, nc7333, 
        nc7334, \A_DOUT_TEMPR95[9] , \A_DOUT_TEMPR95[8] , 
        \A_DOUT_TEMPR95[7] , \A_DOUT_TEMPR95[6] , \A_DOUT_TEMPR95[5] })
        , .B_DOUT({nc7335, nc7336, nc7337, nc7338, nc7339, nc7340, 
        nc7341, nc7342, nc7343, nc7344, nc7345, nc7346, nc7347, nc7348, 
        nc7349, \B_DOUT_TEMPR95[9] , \B_DOUT_TEMPR95[8] , 
        \B_DOUT_TEMPR95[7] , \B_DOUT_TEMPR95[6] , \B_DOUT_TEMPR95[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[95][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2893 (.A(\B_DOUT_TEMPR95[20] ), .B(\B_DOUT_TEMPR96[20] ), 
        .C(\B_DOUT_TEMPR97[20] ), .D(\B_DOUT_TEMPR98[20] ), .Y(
        OR4_2893_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%44%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R44C2 (
        .A_DOUT({nc7350, nc7351, nc7352, nc7353, nc7354, nc7355, 
        nc7356, nc7357, nc7358, nc7359, nc7360, nc7361, nc7362, nc7363, 
        nc7364, \A_DOUT_TEMPR44[14] , \A_DOUT_TEMPR44[13] , 
        \A_DOUT_TEMPR44[12] , \A_DOUT_TEMPR44[11] , 
        \A_DOUT_TEMPR44[10] }), .B_DOUT({nc7365, nc7366, nc7367, 
        nc7368, nc7369, nc7370, nc7371, nc7372, nc7373, nc7374, nc7375, 
        nc7376, nc7377, nc7378, nc7379, \B_DOUT_TEMPR44[14] , 
        \B_DOUT_TEMPR44[13] , \B_DOUT_TEMPR44[12] , 
        \B_DOUT_TEMPR44[11] , \B_DOUT_TEMPR44[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[44][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENB[14]  (.A(B_WBYTE_EN[7]), .B(
        B_WEN), .Y(\WBYTEENB[14] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%85%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R85C6 (
        .A_DOUT({nc7380, nc7381, nc7382, nc7383, nc7384, nc7385, 
        nc7386, nc7387, nc7388, nc7389, nc7390, nc7391, nc7392, nc7393, 
        nc7394, \A_DOUT_TEMPR85[34] , \A_DOUT_TEMPR85[33] , 
        \A_DOUT_TEMPR85[32] , \A_DOUT_TEMPR85[31] , 
        \A_DOUT_TEMPR85[30] }), .B_DOUT({nc7395, nc7396, nc7397, 
        nc7398, nc7399, nc7400, nc7401, nc7402, nc7403, nc7404, nc7405, 
        nc7406, nc7407, nc7408, nc7409, \B_DOUT_TEMPR85[34] , 
        \B_DOUT_TEMPR85[33] , \B_DOUT_TEMPR85[32] , 
        \B_DOUT_TEMPR85[31] , \B_DOUT_TEMPR85[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[85][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%105%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R105C3 (
        .A_DOUT({nc7410, nc7411, nc7412, nc7413, nc7414, nc7415, 
        nc7416, nc7417, nc7418, nc7419, nc7420, nc7421, nc7422, nc7423, 
        nc7424, \A_DOUT_TEMPR105[19] , \A_DOUT_TEMPR105[18] , 
        \A_DOUT_TEMPR105[17] , \A_DOUT_TEMPR105[16] , 
        \A_DOUT_TEMPR105[15] }), .B_DOUT({nc7425, nc7426, nc7427, 
        nc7428, nc7429, nc7430, nc7431, nc7432, nc7433, nc7434, nc7435, 
        nc7436, nc7437, nc7438, nc7439, \B_DOUT_TEMPR105[19] , 
        \B_DOUT_TEMPR105[18] , \B_DOUT_TEMPR105[17] , 
        \B_DOUT_TEMPR105[16] , \B_DOUT_TEMPR105[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[105][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2317 (.A(\A_DOUT_TEMPR95[8] ), .B(\A_DOUT_TEMPR96[8] ), .C(
        \A_DOUT_TEMPR97[8] ), .D(\A_DOUT_TEMPR98[8] ), .Y(OR4_2317_Y));
    OR4 OR4_2212 (.A(OR4_1540_Y), .B(OR4_1988_Y), .C(OR4_2630_Y), .D(
        OR4_1801_Y), .Y(OR4_2212_Y));
    OR4 OR4_1916 (.A(\B_DOUT_TEMPR75[15] ), .B(\B_DOUT_TEMPR76[15] ), 
        .C(\B_DOUT_TEMPR77[15] ), .D(\B_DOUT_TEMPR78[15] ), .Y(
        OR4_1916_Y));
    OR4 OR4_2188 (.A(\A_DOUT_TEMPR40[23] ), .B(\A_DOUT_TEMPR41[23] ), 
        .C(\A_DOUT_TEMPR42[23] ), .D(\A_DOUT_TEMPR43[23] ), .Y(
        OR4_2188_Y));
    OR4 OR4_2799 (.A(\B_DOUT_TEMPR20[4] ), .B(\B_DOUT_TEMPR21[4] ), .C(
        \B_DOUT_TEMPR22[4] ), .D(\B_DOUT_TEMPR23[4] ), .Y(OR4_2799_Y));
    OR4 OR4_1643 (.A(\A_DOUT_TEMPR91[27] ), .B(\A_DOUT_TEMPR92[27] ), 
        .C(\A_DOUT_TEMPR93[27] ), .D(\A_DOUT_TEMPR94[27] ), .Y(
        OR4_1643_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%58%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R58C0 (
        .A_DOUT({nc7440, nc7441, nc7442, nc7443, nc7444, nc7445, 
        nc7446, nc7447, nc7448, nc7449, nc7450, nc7451, nc7452, nc7453, 
        nc7454, \A_DOUT_TEMPR58[4] , \A_DOUT_TEMPR58[3] , 
        \A_DOUT_TEMPR58[2] , \A_DOUT_TEMPR58[1] , \A_DOUT_TEMPR58[0] })
        , .B_DOUT({nc7455, nc7456, nc7457, nc7458, nc7459, nc7460, 
        nc7461, nc7462, nc7463, nc7464, nc7465, nc7466, nc7467, nc7468, 
        nc7469, \B_DOUT_TEMPR58[4] , \B_DOUT_TEMPR58[3] , 
        \B_DOUT_TEMPR58[2] , \B_DOUT_TEMPR58[1] , \B_DOUT_TEMPR58[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[58][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2632 (.A(\A_DOUT_TEMPR16[10] ), .B(\A_DOUT_TEMPR17[10] ), 
        .C(\A_DOUT_TEMPR18[10] ), .D(\A_DOUT_TEMPR19[10] ), .Y(
        OR4_2632_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%11%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R11C3 (
        .A_DOUT({nc7470, nc7471, nc7472, nc7473, nc7474, nc7475, 
        nc7476, nc7477, nc7478, nc7479, nc7480, nc7481, nc7482, nc7483, 
        nc7484, \A_DOUT_TEMPR11[19] , \A_DOUT_TEMPR11[18] , 
        \A_DOUT_TEMPR11[17] , \A_DOUT_TEMPR11[16] , 
        \A_DOUT_TEMPR11[15] }), .B_DOUT({nc7485, nc7486, nc7487, 
        nc7488, nc7489, nc7490, nc7491, nc7492, nc7493, nc7494, nc7495, 
        nc7496, nc7497, nc7498, nc7499, \B_DOUT_TEMPR11[19] , 
        \B_DOUT_TEMPR11[18] , \B_DOUT_TEMPR11[17] , 
        \B_DOUT_TEMPR11[16] , \B_DOUT_TEMPR11[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[11][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[37]  (.A(OR4_1575_Y), .B(OR4_297_Y), .C(OR4_2318_Y)
        , .D(OR4_480_Y), .Y(A_DOUT[37]));
    OR4 OR4_13 (.A(OR4_568_Y), .B(OR4_379_Y), .C(OR2_7_Y), .D(
        \B_DOUT_TEMPR74[34] ), .Y(OR4_13_Y));
    OR4 OR4_739 (.A(\A_DOUT_TEMPR60[8] ), .B(\A_DOUT_TEMPR61[8] ), .C(
        \A_DOUT_TEMPR62[8] ), .D(\A_DOUT_TEMPR63[8] ), .Y(OR4_739_Y));
    OR4 OR4_1949 (.A(\A_DOUT_TEMPR99[32] ), .B(\A_DOUT_TEMPR100[32] ), 
        .C(\A_DOUT_TEMPR101[32] ), .D(\A_DOUT_TEMPR102[32] ), .Y(
        OR4_1949_Y));
    OR4 OR4_662 (.A(\A_DOUT_TEMPR40[8] ), .B(\A_DOUT_TEMPR41[8] ), .C(
        \A_DOUT_TEMPR42[8] ), .D(\A_DOUT_TEMPR43[8] ), .Y(OR4_662_Y));
    OR4 OR4_486 (.A(OR4_2081_Y), .B(OR4_2837_Y), .C(OR4_2351_Y), .D(
        OR4_1315_Y), .Y(OR4_486_Y));
    OR4 OR4_1632 (.A(\A_DOUT_TEMPR75[22] ), .B(\A_DOUT_TEMPR76[22] ), 
        .C(\A_DOUT_TEMPR77[22] ), .D(\A_DOUT_TEMPR78[22] ), .Y(
        OR4_1632_Y));
    OR4 OR4_1381 (.A(OR4_1858_Y), .B(OR4_69_Y), .C(OR4_757_Y), .D(
        OR4_1083_Y), .Y(OR4_1381_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%117%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R117C3 (
        .A_DOUT({nc7500, nc7501, nc7502, nc7503, nc7504, nc7505, 
        nc7506, nc7507, nc7508, nc7509, nc7510, nc7511, nc7512, nc7513, 
        nc7514, \A_DOUT_TEMPR117[19] , \A_DOUT_TEMPR117[18] , 
        \A_DOUT_TEMPR117[17] , \A_DOUT_TEMPR117[16] , 
        \A_DOUT_TEMPR117[15] }), .B_DOUT({nc7515, nc7516, nc7517, 
        nc7518, nc7519, nc7520, nc7521, nc7522, nc7523, nc7524, nc7525, 
        nc7526, nc7527, nc7528, nc7529, \B_DOUT_TEMPR117[19] , 
        \B_DOUT_TEMPR117[18] , \B_DOUT_TEMPR117[17] , 
        \B_DOUT_TEMPR117[16] , \B_DOUT_TEMPR117[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[117][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2932 (.A(OR4_1937_Y), .B(OR4_884_Y), .C(OR4_2529_Y), .D(
        OR4_477_Y), .Y(OR4_2932_Y));
    OR4 OR4_635 (.A(\B_DOUT_TEMPR28[38] ), .B(\B_DOUT_TEMPR29[38] ), 
        .C(\B_DOUT_TEMPR30[38] ), .D(\B_DOUT_TEMPR31[38] ), .Y(
        OR4_635_Y));
    OR4 OR4_904 (.A(\A_DOUT_TEMPR28[22] ), .B(\A_DOUT_TEMPR29[22] ), 
        .C(\A_DOUT_TEMPR30[22] ), .D(\A_DOUT_TEMPR31[22] ), .Y(
        OR4_904_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%43%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R43C7 (
        .A_DOUT({nc7530, nc7531, nc7532, nc7533, nc7534, nc7535, 
        nc7536, nc7537, nc7538, nc7539, nc7540, nc7541, nc7542, nc7543, 
        nc7544, \A_DOUT_TEMPR43[39] , \A_DOUT_TEMPR43[38] , 
        \A_DOUT_TEMPR43[37] , \A_DOUT_TEMPR43[36] , 
        \A_DOUT_TEMPR43[35] }), .B_DOUT({nc7545, nc7546, nc7547, 
        nc7548, nc7549, nc7550, nc7551, nc7552, nc7553, nc7554, nc7555, 
        nc7556, nc7557, nc7558, nc7559, \B_DOUT_TEMPR43[39] , 
        \B_DOUT_TEMPR43[38] , \B_DOUT_TEMPR43[37] , 
        \B_DOUT_TEMPR43[36] , \B_DOUT_TEMPR43[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[43][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1881 (.A(\A_DOUT_TEMPR75[23] ), .B(\A_DOUT_TEMPR76[23] ), 
        .C(\A_DOUT_TEMPR77[23] ), .D(\A_DOUT_TEMPR78[23] ), .Y(
        OR4_1881_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%64%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R64C6 (
        .A_DOUT({nc7560, nc7561, nc7562, nc7563, nc7564, nc7565, 
        nc7566, nc7567, nc7568, nc7569, nc7570, nc7571, nc7572, nc7573, 
        nc7574, \A_DOUT_TEMPR64[34] , \A_DOUT_TEMPR64[33] , 
        \A_DOUT_TEMPR64[32] , \A_DOUT_TEMPR64[31] , 
        \A_DOUT_TEMPR64[30] }), .B_DOUT({nc7575, nc7576, nc7577, 
        nc7578, nc7579, nc7580, nc7581, nc7582, nc7583, nc7584, nc7585, 
        nc7586, nc7587, nc7588, nc7589, \B_DOUT_TEMPR64[34] , 
        \B_DOUT_TEMPR64[33] , \B_DOUT_TEMPR64[32] , 
        \B_DOUT_TEMPR64[31] , \B_DOUT_TEMPR64[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[64][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_150 (.A(\A_DOUT_TEMPR111[37] ), .B(\A_DOUT_TEMPR112[37] ), 
        .C(\A_DOUT_TEMPR113[37] ), .D(\A_DOUT_TEMPR114[37] ), .Y(
        OR4_150_Y));
    OR4 OR4_2196 (.A(OR4_965_Y), .B(OR4_1852_Y), .C(OR4_1497_Y), .D(
        OR4_3011_Y), .Y(OR4_2196_Y));
    OR4 OR4_2883 (.A(\A_DOUT_TEMPR95[7] ), .B(\A_DOUT_TEMPR96[7] ), .C(
        \A_DOUT_TEMPR97[7] ), .D(\A_DOUT_TEMPR98[7] ), .Y(OR4_2883_Y));
    OR4 OR4_2954 (.A(\A_DOUT_TEMPR32[29] ), .B(\A_DOUT_TEMPR33[29] ), 
        .C(\A_DOUT_TEMPR34[29] ), .D(\A_DOUT_TEMPR35[29] ), .Y(
        OR4_2954_Y));
    OR4 OR4_2598 (.A(\B_DOUT_TEMPR64[24] ), .B(\B_DOUT_TEMPR65[24] ), 
        .C(\B_DOUT_TEMPR66[24] ), .D(\B_DOUT_TEMPR67[24] ), .Y(
        OR4_2598_Y));
    OR4 OR4_2414 (.A(\B_DOUT_TEMPR44[39] ), .B(\B_DOUT_TEMPR45[39] ), 
        .C(\B_DOUT_TEMPR46[39] ), .D(\B_DOUT_TEMPR47[39] ), .Y(
        OR4_2414_Y));
    OR4 OR4_1932 (.A(\A_DOUT_TEMPR83[8] ), .B(\A_DOUT_TEMPR84[8] ), .C(
        \A_DOUT_TEMPR85[8] ), .D(\A_DOUT_TEMPR86[8] ), .Y(OR4_1932_Y));
    OR4 OR4_239 (.A(\A_DOUT_TEMPR79[34] ), .B(\A_DOUT_TEMPR80[34] ), 
        .C(\A_DOUT_TEMPR81[34] ), .D(\A_DOUT_TEMPR82[34] ), .Y(
        OR4_239_Y));
    OR4 OR4_92 (.A(\B_DOUT_TEMPR64[20] ), .B(\B_DOUT_TEMPR65[20] ), .C(
        \B_DOUT_TEMPR66[20] ), .D(\B_DOUT_TEMPR67[20] ), .Y(OR4_92_Y));
    OR4 OR4_2572 (.A(\A_DOUT_TEMPR75[27] ), .B(\A_DOUT_TEMPR76[27] ), 
        .C(\A_DOUT_TEMPR77[27] ), .D(\A_DOUT_TEMPR78[27] ), .Y(
        OR4_2572_Y));
    OR4 OR4_2956 (.A(\B_DOUT_TEMPR48[36] ), .B(\B_DOUT_TEMPR49[36] ), 
        .C(\B_DOUT_TEMPR50[36] ), .D(\B_DOUT_TEMPR51[36] ), .Y(
        OR4_2956_Y));
    OR4 OR4_2789 (.A(\B_DOUT_TEMPR0[10] ), .B(\B_DOUT_TEMPR1[10] ), .C(
        \B_DOUT_TEMPR2[10] ), .D(\B_DOUT_TEMPR3[10] ), .Y(OR4_2789_Y));
    OR4 OR4_2923 (.A(\B_DOUT_TEMPR95[16] ), .B(\B_DOUT_TEMPR96[16] ), 
        .C(\B_DOUT_TEMPR97[16] ), .D(\B_DOUT_TEMPR98[16] ), .Y(
        OR4_2923_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[22]  (.A(CFG3_0_Y), .B(CFG3_3_Y)
        , .Y(\BLKX2[22] ));
    OR4 OR4_733 (.A(OR4_862_Y), .B(OR4_1655_Y), .C(OR2_24_Y), .D(
        \A_DOUT_TEMPR74[25] ), .Y(OR4_733_Y));
    OR4 OR4_1744 (.A(\B_DOUT_TEMPR83[36] ), .B(\B_DOUT_TEMPR84[36] ), 
        .C(\B_DOUT_TEMPR85[36] ), .D(\B_DOUT_TEMPR86[36] ), .Y(
        OR4_1744_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[21]  (.A(CFG3_1_Y), .B(CFG3_3_Y)
        , .Y(\BLKX2[21] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%106%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R106C3 (
        .A_DOUT({nc7590, nc7591, nc7592, nc7593, nc7594, nc7595, 
        nc7596, nc7597, nc7598, nc7599, nc7600, nc7601, nc7602, nc7603, 
        nc7604, \A_DOUT_TEMPR106[19] , \A_DOUT_TEMPR106[18] , 
        \A_DOUT_TEMPR106[17] , \A_DOUT_TEMPR106[16] , 
        \A_DOUT_TEMPR106[15] }), .B_DOUT({nc7605, nc7606, nc7607, 
        nc7608, nc7609, nc7610, nc7611, nc7612, nc7613, nc7614, nc7615, 
        nc7616, nc7617, nc7618, nc7619, \B_DOUT_TEMPR106[19] , 
        \B_DOUT_TEMPR106[18] , \B_DOUT_TEMPR106[17] , 
        \B_DOUT_TEMPR106[16] , \B_DOUT_TEMPR106[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[106][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_658 (.A(\B_DOUT_TEMPR107[3] ), .B(\B_DOUT_TEMPR108[3] ), 
        .C(\B_DOUT_TEMPR109[3] ), .D(\B_DOUT_TEMPR110[3] ), .Y(
        OR4_658_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%23%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R23C5 (
        .A_DOUT({nc7620, nc7621, nc7622, nc7623, nc7624, nc7625, 
        nc7626, nc7627, nc7628, nc7629, nc7630, nc7631, nc7632, nc7633, 
        nc7634, \A_DOUT_TEMPR23[29] , \A_DOUT_TEMPR23[28] , 
        \A_DOUT_TEMPR23[27] , \A_DOUT_TEMPR23[26] , 
        \A_DOUT_TEMPR23[25] }), .B_DOUT({nc7635, nc7636, nc7637, 
        nc7638, nc7639, nc7640, nc7641, nc7642, nc7643, nc7644, nc7645, 
        nc7646, nc7647, nc7648, nc7649, \B_DOUT_TEMPR23[29] , 
        \B_DOUT_TEMPR23[28] , \B_DOUT_TEMPR23[27] , 
        \B_DOUT_TEMPR23[26] , \B_DOUT_TEMPR23[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[23][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR2 OR2_77 (.A(\A_DOUT_TEMPR72[2] ), .B(\A_DOUT_TEMPR73[2] ), .Y(
        OR2_77_Y));
    OR4 OR4_0 (.A(\B_DOUT_TEMPR60[34] ), .B(\B_DOUT_TEMPR61[34] ), .C(
        \B_DOUT_TEMPR62[34] ), .D(\B_DOUT_TEMPR63[34] ), .Y(OR4_0_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%10%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R10C2 (
        .A_DOUT({nc7650, nc7651, nc7652, nc7653, nc7654, nc7655, 
        nc7656, nc7657, nc7658, nc7659, nc7660, nc7661, nc7662, nc7663, 
        nc7664, \A_DOUT_TEMPR10[14] , \A_DOUT_TEMPR10[13] , 
        \A_DOUT_TEMPR10[12] , \A_DOUT_TEMPR10[11] , 
        \A_DOUT_TEMPR10[10] }), .B_DOUT({nc7665, nc7666, nc7667, 
        nc7668, nc7669, nc7670, nc7671, nc7672, nc7673, nc7674, nc7675, 
        nc7676, nc7677, nc7678, nc7679, \B_DOUT_TEMPR10[14] , 
        \B_DOUT_TEMPR10[13] , \B_DOUT_TEMPR10[12] , 
        \B_DOUT_TEMPR10[11] , \B_DOUT_TEMPR10[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[10][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1441 (.A(\A_DOUT_TEMPR95[16] ), .B(\A_DOUT_TEMPR96[16] ), 
        .C(\A_DOUT_TEMPR97[16] ), .D(\A_DOUT_TEMPR98[16] ), .Y(
        OR4_1441_Y));
    OR4 OR4_1178 (.A(\B_DOUT_TEMPR52[33] ), .B(\B_DOUT_TEMPR53[33] ), 
        .C(\B_DOUT_TEMPR54[33] ), .D(\B_DOUT_TEMPR55[33] ), .Y(
        OR4_1178_Y));
    OR4 OR4_2149 (.A(\A_DOUT_TEMPR52[26] ), .B(\A_DOUT_TEMPR53[26] ), 
        .C(\A_DOUT_TEMPR54[26] ), .D(\A_DOUT_TEMPR55[26] ), .Y(
        OR4_2149_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%97%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R97C5 (
        .A_DOUT({nc7680, nc7681, nc7682, nc7683, nc7684, nc7685, 
        nc7686, nc7687, nc7688, nc7689, nc7690, nc7691, nc7692, nc7693, 
        nc7694, \A_DOUT_TEMPR97[29] , \A_DOUT_TEMPR97[28] , 
        \A_DOUT_TEMPR97[27] , \A_DOUT_TEMPR97[26] , 
        \A_DOUT_TEMPR97[25] }), .B_DOUT({nc7695, nc7696, nc7697, 
        nc7698, nc7699, nc7700, nc7701, nc7702, nc7703, nc7704, nc7705, 
        nc7706, nc7707, nc7708, nc7709, \B_DOUT_TEMPR97[29] , 
        \B_DOUT_TEMPR97[28] , \B_DOUT_TEMPR97[27] , 
        \B_DOUT_TEMPR97[26] , \B_DOUT_TEMPR97[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[97][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2186 (.A(\B_DOUT_TEMPR16[15] ), .B(\B_DOUT_TEMPR17[15] ), 
        .C(\B_DOUT_TEMPR18[15] ), .D(\B_DOUT_TEMPR19[15] ), .Y(
        OR4_2186_Y));
    OR4 OR4_1868 (.A(\A_DOUT_TEMPR36[21] ), .B(\A_DOUT_TEMPR37[21] ), 
        .C(\A_DOUT_TEMPR38[21] ), .D(\A_DOUT_TEMPR39[21] ), .Y(
        OR4_1868_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[23]  (.A(CFG3_2_Y), .B(
        CFG3_21_Y), .Y(\BLKY2[23] ));
    OR4 OR4_2588 (.A(OR4_627_Y), .B(OR4_2708_Y), .C(OR4_2923_Y), .D(
        OR4_2723_Y), .Y(OR4_2588_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%55%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R55C0 (
        .A_DOUT({nc7710, nc7711, nc7712, nc7713, nc7714, nc7715, 
        nc7716, nc7717, nc7718, nc7719, nc7720, nc7721, nc7722, nc7723, 
        nc7724, \A_DOUT_TEMPR55[4] , \A_DOUT_TEMPR55[3] , 
        \A_DOUT_TEMPR55[2] , \A_DOUT_TEMPR55[1] , \A_DOUT_TEMPR55[0] })
        , .B_DOUT({nc7725, nc7726, nc7727, nc7728, nc7729, nc7730, 
        nc7731, nc7732, nc7733, nc7734, nc7735, nc7736, nc7737, nc7738, 
        nc7739, \B_DOUT_TEMPR55[4] , \B_DOUT_TEMPR55[3] , 
        \B_DOUT_TEMPR55[2] , \B_DOUT_TEMPR55[1] , \B_DOUT_TEMPR55[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[55][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1552 (.A(OR4_1893_Y), .B(OR4_2171_Y), .C(OR4_751_Y), .D(
        OR4_1665_Y), .Y(OR4_1552_Y));
    OR4 OR4_238 (.A(OR4_2066_Y), .B(OR4_584_Y), .C(OR4_1416_Y), .D(
        OR4_431_Y), .Y(OR4_238_Y));
    OR4 OR4_312 (.A(\A_DOUT_TEMPR52[0] ), .B(\A_DOUT_TEMPR53[0] ), .C(
        \A_DOUT_TEMPR54[0] ), .D(\A_DOUT_TEMPR55[0] ), .Y(OR4_312_Y));
    OR4 OR4_2321 (.A(\B_DOUT_TEMPR28[21] ), .B(\B_DOUT_TEMPR29[21] ), 
        .C(\B_DOUT_TEMPR30[21] ), .D(\B_DOUT_TEMPR31[21] ), .Y(
        OR4_2321_Y));
    OR4 OR4_951 (.A(\A_DOUT_TEMPR12[25] ), .B(\A_DOUT_TEMPR13[25] ), 
        .C(\A_DOUT_TEMPR14[25] ), .D(\A_DOUT_TEMPR15[25] ), .Y(
        OR4_951_Y));
    OR4 OR4_1873 (.A(\A_DOUT_TEMPR48[17] ), .B(\A_DOUT_TEMPR49[17] ), 
        .C(\A_DOUT_TEMPR50[17] ), .D(\A_DOUT_TEMPR51[17] ), .Y(
        OR4_1873_Y));
    OR4 OR4_2821 (.A(OR4_1866_Y), .B(OR4_116_Y), .C(OR4_2898_Y), .D(
        OR4_452_Y), .Y(OR4_2821_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%38%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R38C0 (
        .A_DOUT({nc7740, nc7741, nc7742, nc7743, nc7744, nc7745, 
        nc7746, nc7747, nc7748, nc7749, nc7750, nc7751, nc7752, nc7753, 
        nc7754, \A_DOUT_TEMPR38[4] , \A_DOUT_TEMPR38[3] , 
        \A_DOUT_TEMPR38[2] , \A_DOUT_TEMPR38[1] , \A_DOUT_TEMPR38[0] })
        , .B_DOUT({nc7755, nc7756, nc7757, nc7758, nc7759, nc7760, 
        nc7761, nc7762, nc7763, nc7764, nc7765, nc7766, nc7767, nc7768, 
        nc7769, \B_DOUT_TEMPR38[4] , \B_DOUT_TEMPR38[3] , 
        \B_DOUT_TEMPR38[2] , \B_DOUT_TEMPR38[1] , \B_DOUT_TEMPR38[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[38][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1779 (.A(\A_DOUT_TEMPR60[12] ), .B(\A_DOUT_TEMPR61[12] ), 
        .C(\A_DOUT_TEMPR62[12] ), .D(\A_DOUT_TEMPR63[12] ), .Y(
        OR4_1779_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%26%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R26C4 (
        .A_DOUT({nc7770, nc7771, nc7772, nc7773, nc7774, nc7775, 
        nc7776, nc7777, nc7778, nc7779, nc7780, nc7781, nc7782, nc7783, 
        nc7784, \A_DOUT_TEMPR26[24] , \A_DOUT_TEMPR26[23] , 
        \A_DOUT_TEMPR26[22] , \A_DOUT_TEMPR26[21] , 
        \A_DOUT_TEMPR26[20] }), .B_DOUT({nc7785, nc7786, nc7787, 
        nc7788, nc7789, nc7790, nc7791, nc7792, nc7793, nc7794, nc7795, 
        nc7796, nc7797, nc7798, nc7799, \B_DOUT_TEMPR26[24] , 
        \B_DOUT_TEMPR26[23] , \B_DOUT_TEMPR26[22] , 
        \B_DOUT_TEMPR26[21] , \B_DOUT_TEMPR26[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[26][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1944 (.A(\A_DOUT_TEMPR79[37] ), .B(\A_DOUT_TEMPR80[37] ), 
        .C(\A_DOUT_TEMPR81[37] ), .D(\A_DOUT_TEMPR82[37] ), .Y(
        OR4_1944_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%43%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R43C0 (
        .A_DOUT({nc7800, nc7801, nc7802, nc7803, nc7804, nc7805, 
        nc7806, nc7807, nc7808, nc7809, nc7810, nc7811, nc7812, nc7813, 
        nc7814, \A_DOUT_TEMPR43[4] , \A_DOUT_TEMPR43[3] , 
        \A_DOUT_TEMPR43[2] , \A_DOUT_TEMPR43[1] , \A_DOUT_TEMPR43[0] })
        , .B_DOUT({nc7815, nc7816, nc7817, nc7818, nc7819, nc7820, 
        nc7821, nc7822, nc7823, nc7824, nc7825, nc7826, nc7827, nc7828, 
        nc7829, \B_DOUT_TEMPR43[4] , \B_DOUT_TEMPR43[3] , 
        \B_DOUT_TEMPR43[2] , \B_DOUT_TEMPR43[1] , \B_DOUT_TEMPR43[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[43][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[3]  (.A(OR4_446_Y), .B(OR4_2276_Y), .C(OR4_867_Y), 
        .D(OR4_222_Y), .Y(A_DOUT[3]));
    OR4 OR4_2439 (.A(\A_DOUT_TEMPR32[30] ), .B(\A_DOUT_TEMPR33[30] ), 
        .C(\A_DOUT_TEMPR34[30] ), .D(\A_DOUT_TEMPR35[30] ), .Y(
        OR4_2439_Y));
    OR4 OR4_2214 (.A(OR4_2620_Y), .B(OR4_390_Y), .C(OR4_2488_Y), .D(
        OR4_1088_Y), .Y(OR4_2214_Y));
    OR4 OR4_1628 (.A(\B_DOUT_TEMPR16[23] ), .B(\B_DOUT_TEMPR17[23] ), 
        .C(\B_DOUT_TEMPR18[23] ), .D(\B_DOUT_TEMPR19[23] ), .Y(
        OR4_1628_Y));
    OR4 OR4_2070 (.A(\B_DOUT_TEMPR12[33] ), .B(\B_DOUT_TEMPR13[33] ), 
        .C(\B_DOUT_TEMPR14[33] ), .D(\B_DOUT_TEMPR15[33] ), .Y(
        OR4_2070_Y));
    OR2 OR2_48 (.A(\A_DOUT_TEMPR72[5] ), .B(\A_DOUT_TEMPR73[5] ), .Y(
        OR2_48_Y));
    OR4 OR4_1946 (.A(OR4_11_Y), .B(OR4_628_Y), .C(OR4_1275_Y), .D(
        OR4_442_Y), .Y(OR4_1946_Y));
    OR4 OR4_479 (.A(\A_DOUT_TEMPR75[29] ), .B(\A_DOUT_TEMPR76[29] ), 
        .C(\A_DOUT_TEMPR77[29] ), .D(\A_DOUT_TEMPR78[29] ), .Y(
        OR4_479_Y));
    OR4 OR4_23 (.A(\B_DOUT_TEMPR68[4] ), .B(\B_DOUT_TEMPR69[4] ), .C(
        \B_DOUT_TEMPR70[4] ), .D(\B_DOUT_TEMPR71[4] ), .Y(OR4_23_Y));
    OR4 OR4_94 (.A(\A_DOUT_TEMPR36[4] ), .B(\A_DOUT_TEMPR37[4] ), .C(
        \A_DOUT_TEMPR38[4] ), .D(\A_DOUT_TEMPR39[4] ), .Y(OR4_94_Y));
    OR2 OR2_70 (.A(\B_DOUT_TEMPR72[21] ), .B(\B_DOUT_TEMPR73[21] ), .Y(
        OR2_70_Y));
    OR4 OR4_1176 (.A(\B_DOUT_TEMPR8[27] ), .B(\B_DOUT_TEMPR9[27] ), .C(
        \B_DOUT_TEMPR10[27] ), .D(\B_DOUT_TEMPR11[27] ), .Y(OR4_1176_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%25%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R25C5 (
        .A_DOUT({nc7830, nc7831, nc7832, nc7833, nc7834, nc7835, 
        nc7836, nc7837, nc7838, nc7839, nc7840, nc7841, nc7842, nc7843, 
        nc7844, \A_DOUT_TEMPR25[29] , \A_DOUT_TEMPR25[28] , 
        \A_DOUT_TEMPR25[27] , \A_DOUT_TEMPR25[26] , 
        \A_DOUT_TEMPR25[25] }), .B_DOUT({nc7845, nc7846, nc7847, 
        nc7848, nc7849, nc7850, nc7851, nc7852, nc7853, nc7854, nc7855, 
        nc7856, nc7857, nc7858, nc7859, \B_DOUT_TEMPR25[29] , 
        \B_DOUT_TEMPR25[28] , \B_DOUT_TEMPR25[27] , 
        \B_DOUT_TEMPR25[26] , \B_DOUT_TEMPR25[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[25][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_629 (.A(\B_DOUT_TEMPR32[18] ), .B(\B_DOUT_TEMPR33[18] ), 
        .C(\B_DOUT_TEMPR34[18] ), .D(\B_DOUT_TEMPR35[18] ), .Y(
        OR4_629_Y));
    OR4 OR4_1439 (.A(\B_DOUT_TEMPR12[3] ), .B(\B_DOUT_TEMPR13[3] ), .C(
        \B_DOUT_TEMPR14[3] ), .D(\B_DOUT_TEMPR15[3] ), .Y(OR4_1439_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%95%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R95C7 (
        .A_DOUT({nc7860, nc7861, nc7862, nc7863, nc7864, nc7865, 
        nc7866, nc7867, nc7868, nc7869, nc7870, nc7871, nc7872, nc7873, 
        nc7874, \A_DOUT_TEMPR95[39] , \A_DOUT_TEMPR95[38] , 
        \A_DOUT_TEMPR95[37] , \A_DOUT_TEMPR95[36] , 
        \A_DOUT_TEMPR95[35] }), .B_DOUT({nc7875, nc7876, nc7877, 
        nc7878, nc7879, nc7880, nc7881, nc7882, nc7883, nc7884, nc7885, 
        nc7886, nc7887, nc7888, nc7889, \B_DOUT_TEMPR95[39] , 
        \B_DOUT_TEMPR95[38] , \B_DOUT_TEMPR95[37] , 
        \B_DOUT_TEMPR95[36] , \B_DOUT_TEMPR95[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[95][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%101%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R101C3 (
        .A_DOUT({nc7890, nc7891, nc7892, nc7893, nc7894, nc7895, 
        nc7896, nc7897, nc7898, nc7899, nc7900, nc7901, nc7902, nc7903, 
        nc7904, \A_DOUT_TEMPR101[19] , \A_DOUT_TEMPR101[18] , 
        \A_DOUT_TEMPR101[17] , \A_DOUT_TEMPR101[16] , 
        \A_DOUT_TEMPR101[15] }), .B_DOUT({nc7905, nc7906, nc7907, 
        nc7908, nc7909, nc7910, nc7911, nc7912, nc7913, nc7914, nc7915, 
        nc7916, nc7917, nc7918, nc7919, \B_DOUT_TEMPR101[19] , 
        \B_DOUT_TEMPR101[18] , \B_DOUT_TEMPR101[17] , 
        \B_DOUT_TEMPR101[16] , \B_DOUT_TEMPR101[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[101][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1578 (.A(\A_DOUT_TEMPR36[23] ), .B(\A_DOUT_TEMPR37[23] ), 
        .C(\A_DOUT_TEMPR38[23] ), .D(\A_DOUT_TEMPR39[23] ), .Y(
        OR4_1578_Y));
    OR4 OR4_137 (.A(\A_DOUT_TEMPR52[35] ), .B(\A_DOUT_TEMPR53[35] ), 
        .C(\A_DOUT_TEMPR54[35] ), .D(\A_DOUT_TEMPR55[35] ), .Y(
        OR4_137_Y));
    OR4 OR4_515 (.A(\A_DOUT_TEMPR107[14] ), .B(\A_DOUT_TEMPR108[14] ), 
        .C(\A_DOUT_TEMPR109[14] ), .D(\A_DOUT_TEMPR110[14] ), .Y(
        OR4_515_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%24%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R24C5 (
        .A_DOUT({nc7920, nc7921, nc7922, nc7923, nc7924, nc7925, 
        nc7926, nc7927, nc7928, nc7929, nc7930, nc7931, nc7932, nc7933, 
        nc7934, \A_DOUT_TEMPR24[29] , \A_DOUT_TEMPR24[28] , 
        \A_DOUT_TEMPR24[27] , \A_DOUT_TEMPR24[26] , 
        \A_DOUT_TEMPR24[25] }), .B_DOUT({nc7935, nc7936, nc7937, 
        nc7938, nc7939, nc7940, nc7941, nc7942, nc7943, nc7944, nc7945, 
        nc7946, nc7947, nc7948, nc7949, \B_DOUT_TEMPR24[29] , 
        \B_DOUT_TEMPR24[28] , \B_DOUT_TEMPR24[27] , 
        \B_DOUT_TEMPR24[26] , \B_DOUT_TEMPR24[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[24][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_3035 (.A(OR4_1257_Y), .B(OR4_2061_Y), .C(OR4_1138_Y), .D(
        OR4_2352_Y), .Y(OR4_3035_Y));
    OR4 OR4_2594 (.A(\A_DOUT_TEMPR115[15] ), .B(\A_DOUT_TEMPR116[15] ), 
        .C(\A_DOUT_TEMPR117[15] ), .D(\A_DOUT_TEMPR118[15] ), .Y(
        OR4_2594_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%47%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R47C7 (
        .A_DOUT({nc7950, nc7951, nc7952, nc7953, nc7954, nc7955, 
        nc7956, nc7957, nc7958, nc7959, nc7960, nc7961, nc7962, nc7963, 
        nc7964, \A_DOUT_TEMPR47[39] , \A_DOUT_TEMPR47[38] , 
        \A_DOUT_TEMPR47[37] , \A_DOUT_TEMPR47[36] , 
        \A_DOUT_TEMPR47[35] }), .B_DOUT({nc7965, nc7966, nc7967, 
        nc7968, nc7969, nc7970, nc7971, nc7972, nc7973, nc7974, nc7975, 
        nc7976, nc7977, nc7978, nc7979, \B_DOUT_TEMPR47[39] , 
        \B_DOUT_TEMPR47[38] , \B_DOUT_TEMPR47[37] , 
        \B_DOUT_TEMPR47[36] , \B_DOUT_TEMPR47[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[47][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2013 (.A(\B_DOUT_TEMPR56[20] ), .B(\B_DOUT_TEMPR57[20] ), 
        .C(\B_DOUT_TEMPR58[20] ), .D(\B_DOUT_TEMPR59[20] ), .Y(
        OR4_2013_Y));
    OR4 OR4_1768 (.A(\A_DOUT_TEMPR52[12] ), .B(\A_DOUT_TEMPR53[12] ), 
        .C(\A_DOUT_TEMPR54[12] ), .D(\A_DOUT_TEMPR55[12] ), .Y(
        OR4_1768_Y));
    OR4 OR4_954 (.A(\A_DOUT_TEMPR87[28] ), .B(\A_DOUT_TEMPR88[28] ), 
        .C(\A_DOUT_TEMPR89[28] ), .D(\A_DOUT_TEMPR90[28] ), .Y(
        OR4_954_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%59%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R59C1 (
        .A_DOUT({nc7980, nc7981, nc7982, nc7983, nc7984, nc7985, 
        nc7986, nc7987, nc7988, nc7989, nc7990, nc7991, nc7992, nc7993, 
        nc7994, \A_DOUT_TEMPR59[9] , \A_DOUT_TEMPR59[8] , 
        \A_DOUT_TEMPR59[7] , \A_DOUT_TEMPR59[6] , \A_DOUT_TEMPR59[5] })
        , .B_DOUT({nc7995, nc7996, nc7997, nc7998, nc7999, nc8000, 
        nc8001, nc8002, nc8003, nc8004, nc8005, nc8006, nc8007, nc8008, 
        nc8009, \B_DOUT_TEMPR59[9] , \B_DOUT_TEMPR59[8] , 
        \B_DOUT_TEMPR59[7] , \B_DOUT_TEMPR59[6] , \B_DOUT_TEMPR59[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[59][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2611 (.A(\A_DOUT_TEMPR75[21] ), .B(\A_DOUT_TEMPR76[21] ), 
        .C(\A_DOUT_TEMPR77[21] ), .D(\A_DOUT_TEMPR78[21] ), .Y(
        OR4_2611_Y));
    OR4 OR4_1050 (.A(OR4_923_Y), .B(OR4_1727_Y), .C(OR4_1411_Y), .D(
        OR4_127_Y), .Y(OR4_1050_Y));
    OR4 OR4_2330 (.A(OR4_1434_Y), .B(OR4_2191_Y), .C(OR4_1406_Y), .D(
        OR4_325_Y), .Y(OR4_2330_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%35%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R35C0 (
        .A_DOUT({nc8010, nc8011, nc8012, nc8013, nc8014, nc8015, 
        nc8016, nc8017, nc8018, nc8019, nc8020, nc8021, nc8022, nc8023, 
        nc8024, \A_DOUT_TEMPR35[4] , \A_DOUT_TEMPR35[3] , 
        \A_DOUT_TEMPR35[2] , \A_DOUT_TEMPR35[1] , \A_DOUT_TEMPR35[0] })
        , .B_DOUT({nc8025, nc8026, nc8027, nc8028, nc8029, nc8030, 
        nc8031, nc8032, nc8033, nc8034, nc8035, nc8036, nc8037, nc8038, 
        nc8039, \B_DOUT_TEMPR35[4] , \B_DOUT_TEMPR35[3] , 
        \B_DOUT_TEMPR35[2] , \B_DOUT_TEMPR35[1] , \B_DOUT_TEMPR35[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[35][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[8] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%76%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R76C0 (
        .A_DOUT({nc8040, nc8041, nc8042, nc8043, nc8044, nc8045, 
        nc8046, nc8047, nc8048, nc8049, nc8050, nc8051, nc8052, nc8053, 
        nc8054, \A_DOUT_TEMPR76[4] , \A_DOUT_TEMPR76[3] , 
        \A_DOUT_TEMPR76[2] , \A_DOUT_TEMPR76[1] , \A_DOUT_TEMPR76[0] })
        , .B_DOUT({nc8055, nc8056, nc8057, nc8058, nc8059, nc8060, 
        nc8061, nc8062, nc8063, nc8064, nc8065, nc8066, nc8067, nc8068, 
        nc8069, \B_DOUT_TEMPR76[4] , \B_DOUT_TEMPR76[3] , 
        \B_DOUT_TEMPR76[2] , \B_DOUT_TEMPR76[1] , \B_DOUT_TEMPR76[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[76][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_923 (.A(OR4_2167_Y), .B(OR4_2477_Y), .C(OR4_1071_Y), .D(
        OR4_1965_Y), .Y(OR4_923_Y));
    OR4 OR4_2437 (.A(\A_DOUT_TEMPR20[15] ), .B(\A_DOUT_TEMPR21[15] ), 
        .C(\A_DOUT_TEMPR22[15] ), .D(\A_DOUT_TEMPR23[15] ), .Y(
        OR4_2437_Y));
    OR4 OR4_2713 (.A(OR4_313_Y), .B(OR4_1408_Y), .C(OR4_3006_Y), .D(
        OR4_372_Y), .Y(OR4_2713_Y));
    OR4 OR4_190 (.A(\A_DOUT_TEMPR107[27] ), .B(\A_DOUT_TEMPR108[27] ), 
        .C(\A_DOUT_TEMPR109[27] ), .D(\A_DOUT_TEMPR110[27] ), .Y(
        OR4_190_Y));
    OR4 OR4_1200 (.A(OR4_1371_Y), .B(OR4_1194_Y), .C(OR4_1135_Y), .D(
        OR4_1885_Y), .Y(OR4_1200_Y));
    OR4 OR4_171 (.A(\B_DOUT_TEMPR79[34] ), .B(\B_DOUT_TEMPR80[34] ), 
        .C(\B_DOUT_TEMPR81[34] ), .D(\B_DOUT_TEMPR82[34] ), .Y(
        OR4_171_Y));
    OR4 OR4_2168 (.A(\B_DOUT_TEMPR16[8] ), .B(\B_DOUT_TEMPR17[8] ), .C(
        \B_DOUT_TEMPR18[8] ), .D(\B_DOUT_TEMPR19[8] ), .Y(OR4_2168_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%85%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R85C2 (
        .A_DOUT({nc8070, nc8071, nc8072, nc8073, nc8074, nc8075, 
        nc8076, nc8077, nc8078, nc8079, nc8080, nc8081, nc8082, nc8083, 
        nc8084, \A_DOUT_TEMPR85[14] , \A_DOUT_TEMPR85[13] , 
        \A_DOUT_TEMPR85[12] , \A_DOUT_TEMPR85[11] , 
        \A_DOUT_TEMPR85[10] }), .B_DOUT({nc8085, nc8086, nc8087, 
        nc8088, nc8089, nc8090, nc8091, nc8092, nc8093, nc8094, nc8095, 
        nc8096, nc8097, nc8098, nc8099, \B_DOUT_TEMPR85[14] , 
        \B_DOUT_TEMPR85[13] , \B_DOUT_TEMPR85[12] , 
        \B_DOUT_TEMPR85[11] , \B_DOUT_TEMPR85[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[85][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1330 (.A(OR4_2895_Y), .B(OR4_2696_Y), .C(OR2_66_Y), .D(
        \A_DOUT_TEMPR74[30] ), .Y(OR4_1330_Y));
    OR4 OR4_1437 (.A(\A_DOUT_TEMPR115[9] ), .B(\A_DOUT_TEMPR116[9] ), 
        .C(\A_DOUT_TEMPR117[9] ), .D(\A_DOUT_TEMPR118[9] ), .Y(
        OR4_1437_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%59%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R59C2 (
        .A_DOUT({nc8100, nc8101, nc8102, nc8103, nc8104, nc8105, 
        nc8106, nc8107, nc8108, nc8109, nc8110, nc8111, nc8112, nc8113, 
        nc8114, \A_DOUT_TEMPR59[14] , \A_DOUT_TEMPR59[13] , 
        \A_DOUT_TEMPR59[12] , \A_DOUT_TEMPR59[11] , 
        \A_DOUT_TEMPR59[10] }), .B_DOUT({nc8115, nc8116, nc8117, 
        nc8118, nc8119, nc8120, nc8121, nc8122, nc8123, nc8124, nc8125, 
        nc8126, nc8127, nc8128, nc8129, \B_DOUT_TEMPR59[14] , 
        \B_DOUT_TEMPR59[13] , \B_DOUT_TEMPR59[12] , 
        \B_DOUT_TEMPR59[11] , \B_DOUT_TEMPR59[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[59][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2115 (.A(\A_DOUT_TEMPR103[16] ), .B(\A_DOUT_TEMPR104[16] ), 
        .C(\A_DOUT_TEMPR105[16] ), .D(\A_DOUT_TEMPR106[16] ), .Y(
        OR4_2115_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%55%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R55C1 (
        .A_DOUT({nc8130, nc8131, nc8132, nc8133, nc8134, nc8135, 
        nc8136, nc8137, nc8138, nc8139, nc8140, nc8141, nc8142, nc8143, 
        nc8144, \A_DOUT_TEMPR55[9] , \A_DOUT_TEMPR55[8] , 
        \A_DOUT_TEMPR55[7] , \A_DOUT_TEMPR55[6] , \A_DOUT_TEMPR55[5] })
        , .B_DOUT({nc8145, nc8146, nc8147, nc8148, nc8149, nc8150, 
        nc8151, nc8152, nc8153, nc8154, nc8155, nc8156, nc8157, nc8158, 
        nc8159, \B_DOUT_TEMPR55[9] , \B_DOUT_TEMPR55[8] , 
        \B_DOUT_TEMPR55[7] , \B_DOUT_TEMPR55[6] , \B_DOUT_TEMPR55[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[55][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2842 (.A(\A_DOUT_TEMPR20[34] ), .B(\A_DOUT_TEMPR21[34] ), 
        .C(\A_DOUT_TEMPR22[34] ), .D(\A_DOUT_TEMPR23[34] ), .Y(
        OR4_2842_Y));
    OR4 OR4_2584 (.A(\B_DOUT_TEMPR111[3] ), .B(\B_DOUT_TEMPR112[3] ), 
        .C(\B_DOUT_TEMPR113[3] ), .D(\B_DOUT_TEMPR114[3] ), .Y(
        OR4_2584_Y));
    OR4 OR4_1987 (.A(\B_DOUT_TEMPR87[23] ), .B(\B_DOUT_TEMPR88[23] ), 
        .C(\B_DOUT_TEMPR89[23] ), .D(\B_DOUT_TEMPR90[23] ), .Y(
        OR4_1987_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%14%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R14C6 (
        .A_DOUT({nc8160, nc8161, nc8162, nc8163, nc8164, nc8165, 
        nc8166, nc8167, nc8168, nc8169, nc8170, nc8171, nc8172, nc8173, 
        nc8174, \A_DOUT_TEMPR14[34] , \A_DOUT_TEMPR14[33] , 
        \A_DOUT_TEMPR14[32] , \A_DOUT_TEMPR14[31] , 
        \A_DOUT_TEMPR14[30] }), .B_DOUT({nc8175, nc8176, nc8177, 
        nc8178, nc8179, nc8180, nc8181, nc8182, nc8183, nc8184, nc8185, 
        nc8186, nc8187, nc8188, nc8189, \B_DOUT_TEMPR14[34] , 
        \B_DOUT_TEMPR14[33] , \B_DOUT_TEMPR14[32] , 
        \B_DOUT_TEMPR14[31] , \B_DOUT_TEMPR14[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[14][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%111%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R111C1 (
        .A_DOUT({nc8190, nc8191, nc8192, nc8193, nc8194, nc8195, 
        nc8196, nc8197, nc8198, nc8199, nc8200, nc8201, nc8202, nc8203, 
        nc8204, \A_DOUT_TEMPR111[9] , \A_DOUT_TEMPR111[8] , 
        \A_DOUT_TEMPR111[7] , \A_DOUT_TEMPR111[6] , 
        \A_DOUT_TEMPR111[5] }), .B_DOUT({nc8205, nc8206, nc8207, 
        nc8208, nc8209, nc8210, nc8211, nc8212, nc8213, nc8214, nc8215, 
        nc8216, nc8217, nc8218, nc8219, \B_DOUT_TEMPR111[9] , 
        \B_DOUT_TEMPR111[8] , \B_DOUT_TEMPR111[7] , 
        \B_DOUT_TEMPR111[6] , \B_DOUT_TEMPR111[5] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[111][1] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[9], 
        B_DIN[8], B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1192 (.A(\B_DOUT_TEMPR32[30] ), .B(\B_DOUT_TEMPR33[30] ), 
        .C(\B_DOUT_TEMPR34[30] ), .D(\B_DOUT_TEMPR35[30] ), .Y(
        OR4_1192_Y));
    OR4 OR4_2476 (.A(\A_DOUT_TEMPR52[37] ), .B(\A_DOUT_TEMPR53[37] ), 
        .C(\A_DOUT_TEMPR54[37] ), .D(\A_DOUT_TEMPR55[37] ), .Y(
        OR4_2476_Y));
    OR4 OR4_2291 (.A(\B_DOUT_TEMPR32[31] ), .B(\B_DOUT_TEMPR33[31] ), 
        .C(\B_DOUT_TEMPR34[31] ), .D(\B_DOUT_TEMPR35[31] ), .Y(
        OR4_2291_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%118%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R118C2 (
        .A_DOUT({nc8220, nc8221, nc8222, nc8223, nc8224, nc8225, 
        nc8226, nc8227, nc8228, nc8229, nc8230, nc8231, nc8232, nc8233, 
        nc8234, \A_DOUT_TEMPR118[14] , \A_DOUT_TEMPR118[13] , 
        \A_DOUT_TEMPR118[12] , \A_DOUT_TEMPR118[11] , 
        \A_DOUT_TEMPR118[10] }), .B_DOUT({nc8235, nc8236, nc8237, 
        nc8238, nc8239, nc8240, nc8241, nc8242, nc8243, nc8244, nc8245, 
        nc8246, nc8247, nc8248, nc8249, \B_DOUT_TEMPR118[14] , 
        \B_DOUT_TEMPR118[13] , \B_DOUT_TEMPR118[12] , 
        \B_DOUT_TEMPR118[11] , \B_DOUT_TEMPR118[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[118][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_409 (.A(\A_DOUT_TEMPR99[3] ), .B(\A_DOUT_TEMPR100[3] ), .C(
        \A_DOUT_TEMPR101[3] ), .D(\A_DOUT_TEMPR102[3] ), .Y(OR4_409_Y));
    OR4 OR4_698 (.A(\A_DOUT_TEMPR68[29] ), .B(\A_DOUT_TEMPR69[29] ), 
        .C(\A_DOUT_TEMPR70[29] ), .D(\A_DOUT_TEMPR71[29] ), .Y(
        OR4_698_Y));
    OR4 OR4_72 (.A(OR4_2427_Y), .B(OR4_1438_Y), .C(OR4_2128_Y), .D(
        OR4_2423_Y), .Y(OR4_72_Y));
    OR4 OR4_2863 (.A(\A_DOUT_TEMPR56[35] ), .B(\A_DOUT_TEMPR57[35] ), 
        .C(\A_DOUT_TEMPR58[35] ), .D(\A_DOUT_TEMPR59[35] ), .Y(
        OR4_2863_Y));
    OR4 OR4_2009 (.A(\B_DOUT_TEMPR12[23] ), .B(\B_DOUT_TEMPR13[23] ), 
        .C(\B_DOUT_TEMPR14[23] ), .D(\B_DOUT_TEMPR15[23] ), .Y(
        OR4_2009_Y));
    OR4 \OR4_B_DOUT[8]  (.A(OR4_2265_Y), .B(OR4_1235_Y), .C(OR4_2700_Y)
        , .D(OR4_2169_Y), .Y(B_DOUT[8]));
    OR4 OR4_2011 (.A(\B_DOUT_TEMPR99[17] ), .B(\B_DOUT_TEMPR100[17] ), 
        .C(\B_DOUT_TEMPR101[17] ), .D(\B_DOUT_TEMPR102[17] ), .Y(
        OR4_2011_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%109%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R109C3 (
        .A_DOUT({nc8250, nc8251, nc8252, nc8253, nc8254, nc8255, 
        nc8256, nc8257, nc8258, nc8259, nc8260, nc8261, nc8262, nc8263, 
        nc8264, \A_DOUT_TEMPR109[19] , \A_DOUT_TEMPR109[18] , 
        \A_DOUT_TEMPR109[17] , \A_DOUT_TEMPR109[16] , 
        \A_DOUT_TEMPR109[15] }), .B_DOUT({nc8265, nc8266, nc8267, 
        nc8268, nc8269, nc8270, nc8271, nc8272, nc8273, nc8274, nc8275, 
        nc8276, nc8277, nc8278, nc8279, \B_DOUT_TEMPR109[19] , 
        \B_DOUT_TEMPR109[18] , \B_DOUT_TEMPR109[17] , 
        \B_DOUT_TEMPR109[16] , \B_DOUT_TEMPR109[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[109][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1306 (.A(\A_DOUT_TEMPR95[19] ), .B(\A_DOUT_TEMPR96[19] ), 
        .C(\A_DOUT_TEMPR97[19] ), .D(\A_DOUT_TEMPR98[19] ), .Y(
        OR4_1306_Y));
    OR4 OR4_2509 (.A(\B_DOUT_TEMPR28[14] ), .B(\B_DOUT_TEMPR29[14] ), 
        .C(\B_DOUT_TEMPR30[14] ), .D(\B_DOUT_TEMPR31[14] ), .Y(
        OR4_2509_Y));
    OR4 OR4_2769 (.A(\B_DOUT_TEMPR36[29] ), .B(\B_DOUT_TEMPR37[29] ), 
        .C(\B_DOUT_TEMPR38[29] ), .D(\B_DOUT_TEMPR39[29] ), .Y(
        OR4_2769_Y));
    OR4 OR4_275 (.A(\A_DOUT_TEMPR60[14] ), .B(\A_DOUT_TEMPR61[14] ), 
        .C(\A_DOUT_TEMPR62[14] ), .D(\A_DOUT_TEMPR63[14] ), .Y(
        OR4_275_Y));
    OR4 OR4_649 (.A(\A_DOUT_TEMPR24[11] ), .B(\A_DOUT_TEMPR25[11] ), 
        .C(\A_DOUT_TEMPR26[11] ), .D(\A_DOUT_TEMPR27[11] ), .Y(
        OR4_649_Y));
    OR4 OR4_2775 (.A(\B_DOUT_TEMPR111[31] ), .B(\B_DOUT_TEMPR112[31] ), 
        .C(\B_DOUT_TEMPR113[31] ), .D(\B_DOUT_TEMPR114[31] ), .Y(
        OR4_2775_Y));
    OR4 OR4_991 (.A(\B_DOUT_TEMPR48[34] ), .B(\B_DOUT_TEMPR49[34] ), 
        .C(\B_DOUT_TEMPR50[34] ), .D(\B_DOUT_TEMPR51[34] ), .Y(
        OR4_991_Y));
    OR4 OR4_1456 (.A(\A_DOUT_TEMPR83[22] ), .B(\A_DOUT_TEMPR84[22] ), 
        .C(\A_DOUT_TEMPR85[22] ), .D(\A_DOUT_TEMPR86[22] ), .Y(
        OR4_1456_Y));
    OR4 OR4_2643 (.A(\B_DOUT_TEMPR40[23] ), .B(\B_DOUT_TEMPR41[23] ), 
        .C(\B_DOUT_TEMPR42[23] ), .D(\B_DOUT_TEMPR43[23] ), .Y(
        OR4_2643_Y));
    OR4 OR4_1880 (.A(OR4_685_Y), .B(OR4_1005_Y), .C(OR4_2600_Y), .D(
        OR4_463_Y), .Y(OR4_1880_Y));
    OR4 OR4_2281 (.A(\A_DOUT_TEMPR111[20] ), .B(\A_DOUT_TEMPR112[20] ), 
        .C(\A_DOUT_TEMPR113[20] ), .D(\A_DOUT_TEMPR114[20] ), .Y(
        OR4_2281_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%74%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R74C2 (
        .A_DOUT({nc8280, nc8281, nc8282, nc8283, nc8284, nc8285, 
        nc8286, nc8287, nc8288, nc8289, nc8290, nc8291, nc8292, nc8293, 
        nc8294, \A_DOUT_TEMPR74[14] , \A_DOUT_TEMPR74[13] , 
        \A_DOUT_TEMPR74[12] , \A_DOUT_TEMPR74[11] , 
        \A_DOUT_TEMPR74[10] }), .B_DOUT({nc8295, nc8296, nc8297, 
        nc8298, nc8299, nc8300, nc8301, nc8302, nc8303, nc8304, nc8305, 
        nc8306, nc8307, nc8308, nc8309, \B_DOUT_TEMPR74[14] , 
        \B_DOUT_TEMPR74[13] , \B_DOUT_TEMPR74[12] , 
        \B_DOUT_TEMPR74[11] , \B_DOUT_TEMPR74[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[74][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2949 (.A(\B_DOUT_TEMPR111[23] ), .B(\B_DOUT_TEMPR112[23] ), 
        .C(\B_DOUT_TEMPR113[23] ), .D(\B_DOUT_TEMPR114[23] ), .Y(
        OR4_2949_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%39%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R39C1 (
        .A_DOUT({nc8310, nc8311, nc8312, nc8313, nc8314, nc8315, 
        nc8316, nc8317, nc8318, nc8319, nc8320, nc8321, nc8322, nc8323, 
        nc8324, \A_DOUT_TEMPR39[9] , \A_DOUT_TEMPR39[8] , 
        \A_DOUT_TEMPR39[7] , \A_DOUT_TEMPR39[6] , \A_DOUT_TEMPR39[5] })
        , .B_DOUT({nc8325, nc8326, nc8327, nc8328, nc8329, nc8330, 
        nc8331, nc8332, nc8333, nc8334, nc8335, nc8336, nc8337, nc8338, 
        nc8339, \B_DOUT_TEMPR39[9] , \B_DOUT_TEMPR39[8] , 
        \B_DOUT_TEMPR39[7] , \B_DOUT_TEMPR39[6] , \B_DOUT_TEMPR39[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[39][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], 
        A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_101 (.A(\B_DOUT_TEMPR64[16] ), .B(\B_DOUT_TEMPR65[16] ), 
        .C(\B_DOUT_TEMPR66[16] ), .D(\B_DOUT_TEMPR67[16] ), .Y(
        OR4_101_Y));
    OR4 OR4_2302 (.A(\A_DOUT_TEMPR12[0] ), .B(\A_DOUT_TEMPR13[0] ), .C(
        \A_DOUT_TEMPR14[0] ), .D(\A_DOUT_TEMPR15[0] ), .Y(OR4_2302_Y));
    OR4 OR4_2166 (.A(\A_DOUT_TEMPR24[37] ), .B(\A_DOUT_TEMPR25[37] ), 
        .C(\A_DOUT_TEMPR26[37] ), .D(\A_DOUT_TEMPR27[37] ), .Y(
        OR4_2166_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%97%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R97C2 (
        .A_DOUT({nc8340, nc8341, nc8342, nc8343, nc8344, nc8345, 
        nc8346, nc8347, nc8348, nc8349, nc8350, nc8351, nc8352, nc8353, 
        nc8354, \A_DOUT_TEMPR97[14] , \A_DOUT_TEMPR97[13] , 
        \A_DOUT_TEMPR97[12] , \A_DOUT_TEMPR97[11] , 
        \A_DOUT_TEMPR97[10] }), .B_DOUT({nc8355, nc8356, nc8357, 
        nc8358, nc8359, nc8360, nc8361, nc8362, nc8363, nc8364, nc8365, 
        nc8366, nc8367, nc8368, nc8369, \B_DOUT_TEMPR97[14] , 
        \B_DOUT_TEMPR97[13] , \B_DOUT_TEMPR97[12] , 
        \B_DOUT_TEMPR97[11] , \B_DOUT_TEMPR97[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[97][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_676 (.A(\A_DOUT_TEMPR56[31] ), .B(\A_DOUT_TEMPR57[31] ), 
        .C(\A_DOUT_TEMPR58[31] ), .D(\A_DOUT_TEMPR59[31] ), .Y(
        OR4_676_Y));
    OR4 OR4_1574 (.A(OR4_2651_Y), .B(OR4_2437_Y), .C(OR4_272_Y), .D(
        OR4_1460_Y), .Y(OR4_1574_Y));
    OR4 OR4_2568 (.A(OR4_952_Y), .B(OR4_1323_Y), .C(OR4_2049_Y), .D(
        OR4_2890_Y), .Y(OR4_2568_Y));
    OR4 OR4_362 (.A(OR4_2635_Y), .B(OR4_2429_Y), .C(OR2_57_Y), .D(
        \B_DOUT_TEMPR74[32] ), .Y(OR4_362_Y));
    OR4 OR4_236 (.A(OR4_723_Y), .B(OR4_2132_Y), .C(OR4_581_Y), .D(
        OR4_2133_Y), .Y(OR4_236_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%28%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R28C4 (
        .A_DOUT({nc8370, nc8371, nc8372, nc8373, nc8374, nc8375, 
        nc8376, nc8377, nc8378, nc8379, nc8380, nc8381, nc8382, nc8383, 
        nc8384, \A_DOUT_TEMPR28[24] , \A_DOUT_TEMPR28[23] , 
        \A_DOUT_TEMPR28[22] , \A_DOUT_TEMPR28[21] , 
        \A_DOUT_TEMPR28[20] }), .B_DOUT({nc8385, nc8386, nc8387, 
        nc8388, nc8389, nc8390, nc8391, nc8392, nc8393, nc8394, nc8395, 
        nc8396, nc8397, nc8398, nc8399, \B_DOUT_TEMPR28[24] , 
        \B_DOUT_TEMPR28[23] , \B_DOUT_TEMPR28[22] , 
        \B_DOUT_TEMPR28[21] , \B_DOUT_TEMPR28[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[28][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2927 (.A(\B_DOUT_TEMPR107[2] ), .B(\B_DOUT_TEMPR108[2] ), 
        .C(\B_DOUT_TEMPR109[2] ), .D(\B_DOUT_TEMPR110[2] ), .Y(
        OR4_2927_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%68%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R68C0 (
        .A_DOUT({nc8400, nc8401, nc8402, nc8403, nc8404, nc8405, 
        nc8406, nc8407, nc8408, nc8409, nc8410, nc8411, nc8412, nc8413, 
        nc8414, \A_DOUT_TEMPR68[4] , \A_DOUT_TEMPR68[3] , 
        \A_DOUT_TEMPR68[2] , \A_DOUT_TEMPR68[1] , \A_DOUT_TEMPR68[0] })
        , .B_DOUT({nc8415, nc8416, nc8417, nc8418, nc8419, nc8420, 
        nc8421, nc8422, nc8423, nc8424, nc8425, nc8426, nc8427, nc8428, 
        nc8429, \B_DOUT_TEMPR68[4] , \B_DOUT_TEMPR68[3] , 
        \B_DOUT_TEMPR68[2] , \B_DOUT_TEMPR68[1] , \B_DOUT_TEMPR68[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[68][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_943 (.A(\B_DOUT_TEMPR68[20] ), .B(\B_DOUT_TEMPR69[20] ), 
        .C(\B_DOUT_TEMPR70[20] ), .D(\B_DOUT_TEMPR71[20] ), .Y(
        OR4_943_Y));
    OR4 OR4_1884 (.A(\B_DOUT_TEMPR0[4] ), .B(\B_DOUT_TEMPR1[4] ), .C(
        \B_DOUT_TEMPR2[4] ), .D(\B_DOUT_TEMPR3[4] ), .Y(OR4_1884_Y));
    OR4 \OR4_B_DOUT[34]  (.A(OR4_2872_Y), .B(OR4_1878_Y), .C(
        OR4_1721_Y), .D(OR4_1510_Y), .Y(B_DOUT[34]));
    OR2 OR2_75 (.A(\B_DOUT_TEMPR72[8] ), .B(\B_DOUT_TEMPR73[8] ), .Y(
        OR2_75_Y));
    OR4 OR4_280 (.A(\A_DOUT_TEMPR20[2] ), .B(\A_DOUT_TEMPR21[2] ), .C(
        \A_DOUT_TEMPR22[2] ), .D(\A_DOUT_TEMPR23[2] ), .Y(OR4_280_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%57%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R57C5 (
        .A_DOUT({nc8430, nc8431, nc8432, nc8433, nc8434, nc8435, 
        nc8436, nc8437, nc8438, nc8439, nc8440, nc8441, nc8442, nc8443, 
        nc8444, \A_DOUT_TEMPR57[29] , \A_DOUT_TEMPR57[28] , 
        \A_DOUT_TEMPR57[27] , \A_DOUT_TEMPR57[26] , 
        \A_DOUT_TEMPR57[25] }), .B_DOUT({nc8445, nc8446, nc8447, 
        nc8448, nc8449, nc8450, nc8451, nc8452, nc8453, nc8454, nc8455, 
        nc8456, nc8457, nc8458, nc8459, \B_DOUT_TEMPR57[29] , 
        \B_DOUT_TEMPR57[28] , \B_DOUT_TEMPR57[27] , 
        \B_DOUT_TEMPR57[26] , \B_DOUT_TEMPR57[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[57][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1755 (.A(OR4_682_Y), .B(OR4_2762_Y), .C(OR4_2969_Y), .D(
        OR4_2783_Y), .Y(OR4_1755_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%39%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R39C2 (
        .A_DOUT({nc8460, nc8461, nc8462, nc8463, nc8464, nc8465, 
        nc8466, nc8467, nc8468, nc8469, nc8470, nc8471, nc8472, nc8473, 
        nc8474, \A_DOUT_TEMPR39[14] , \A_DOUT_TEMPR39[13] , 
        \A_DOUT_TEMPR39[12] , \A_DOUT_TEMPR39[11] , 
        \A_DOUT_TEMPR39[10] }), .B_DOUT({nc8475, nc8476, nc8477, 
        nc8478, nc8479, nc8480, nc8481, nc8482, nc8483, nc8484, nc8485, 
        nc8486, nc8487, nc8488, nc8489, \B_DOUT_TEMPR39[14] , 
        \B_DOUT_TEMPR39[13] , \B_DOUT_TEMPR39[12] , 
        \B_DOUT_TEMPR39[11] , \B_DOUT_TEMPR39[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[39][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%35%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R35C1 (
        .A_DOUT({nc8490, nc8491, nc8492, nc8493, nc8494, nc8495, 
        nc8496, nc8497, nc8498, nc8499, nc8500, nc8501, nc8502, nc8503, 
        nc8504, \A_DOUT_TEMPR35[9] , \A_DOUT_TEMPR35[8] , 
        \A_DOUT_TEMPR35[7] , \A_DOUT_TEMPR35[6] , \A_DOUT_TEMPR35[5] })
        , .B_DOUT({nc8505, nc8506, nc8507, nc8508, nc8509, nc8510, 
        nc8511, nc8512, nc8513, nc8514, nc8515, nc8516, nc8517, nc8518, 
        nc8519, \B_DOUT_TEMPR35[9] , \B_DOUT_TEMPR35[8] , 
        \B_DOUT_TEMPR35[7] , \B_DOUT_TEMPR35[6] , \B_DOUT_TEMPR35[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[35][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[8] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], 
        A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1829 (.A(\B_DOUT_TEMPR4[3] ), .B(\B_DOUT_TEMPR5[3] ), .C(
        \B_DOUT_TEMPR6[3] ), .D(\B_DOUT_TEMPR7[3] ), .Y(OR4_1829_Y));
    OR4 OR4_680 (.A(OR4_2029_Y), .B(OR4_1234_Y), .C(OR4_169_Y), .D(
        OR4_491_Y), .Y(OR4_680_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%73%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R73C7 (
        .A_DOUT({nc8520, nc8521, nc8522, nc8523, nc8524, nc8525, 
        nc8526, nc8527, nc8528, nc8529, nc8530, nc8531, nc8532, nc8533, 
        nc8534, \A_DOUT_TEMPR73[39] , \A_DOUT_TEMPR73[38] , 
        \A_DOUT_TEMPR73[37] , \A_DOUT_TEMPR73[36] , 
        \A_DOUT_TEMPR73[35] }), .B_DOUT({nc8535, nc8536, nc8537, 
        nc8538, nc8539, nc8540, nc8541, nc8542, nc8543, nc8544, nc8545, 
        nc8546, nc8547, nc8548, nc8549, \B_DOUT_TEMPR73[39] , 
        \B_DOUT_TEMPR73[38] , \B_DOUT_TEMPR73[37] , 
        \B_DOUT_TEMPR73[36] , \B_DOUT_TEMPR73[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[73][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2744 (.A(OR4_2055_Y), .B(OR4_20_Y), .C(OR4_688_Y), .D(
        OR4_2340_Y), .Y(OR4_2744_Y));
    OR4 OR4_2441 (.A(\A_DOUT_TEMPR0[12] ), .B(\A_DOUT_TEMPR1[12] ), .C(
        \A_DOUT_TEMPR2[12] ), .D(\A_DOUT_TEMPR3[12] ), .Y(OR4_2441_Y));
    OR4 OR4_205 (.A(\A_DOUT_TEMPR12[7] ), .B(\A_DOUT_TEMPR13[7] ), .C(
        \A_DOUT_TEMPR14[7] ), .D(\A_DOUT_TEMPR15[7] ), .Y(OR4_205_Y));
    OR4 OR4_74 (.A(\B_DOUT_TEMPR115[35] ), .B(\B_DOUT_TEMPR116[35] ), 
        .C(\B_DOUT_TEMPR117[35] ), .D(\B_DOUT_TEMPR118[35] ), .Y(
        OR4_74_Y));
    OR4 OR4_1121 (.A(\A_DOUT_TEMPR20[9] ), .B(\A_DOUT_TEMPR21[9] ), .C(
        \A_DOUT_TEMPR22[9] ), .D(\A_DOUT_TEMPR23[9] ), .Y(OR4_1121_Y));
    OR4 OR4_994 (.A(\A_DOUT_TEMPR24[14] ), .B(\A_DOUT_TEMPR25[14] ), 
        .C(\A_DOUT_TEMPR26[14] ), .D(\A_DOUT_TEMPR27[14] ), .Y(
        OR4_994_Y));
    OR4 OR4_2505 (.A(OR4_786_Y), .B(OR4_1112_Y), .C(OR4_719_Y), .D(
        OR4_1133_Y), .Y(OR4_2505_Y));
    OR4 OR4_1402 (.A(OR4_1823_Y), .B(OR4_871_Y), .C(OR4_1081_Y), .D(
        OR4_881_Y), .Y(OR4_1402_Y));
    OR4 OR4_2820 (.A(OR4_1246_Y), .B(OR4_2158_Y), .C(OR4_1342_Y), .D(
        OR4_1649_Y), .Y(OR4_2820_Y));
    OR4 OR4_1271 (.A(\A_DOUT_TEMPR79[33] ), .B(\A_DOUT_TEMPR80[33] ), 
        .C(\A_DOUT_TEMPR81[33] ), .D(\A_DOUT_TEMPR82[33] ), .Y(
        OR4_1271_Y));
    OR4 OR4_174 (.A(\B_DOUT_TEMPR56[2] ), .B(\B_DOUT_TEMPR57[2] ), .C(
        \B_DOUT_TEMPR58[2] ), .D(\B_DOUT_TEMPR59[2] ), .Y(OR4_174_Y));
    OR4 OR4_374 (.A(OR4_1542_Y), .B(OR4_1846_Y), .C(OR4_1479_Y), .D(
        OR4_1870_Y), .Y(OR4_374_Y));
    OR4 OR4_565 (.A(\B_DOUT_TEMPR103[11] ), .B(\B_DOUT_TEMPR104[11] ), 
        .C(\B_DOUT_TEMPR105[11] ), .D(\B_DOUT_TEMPR106[11] ), .Y(
        OR4_565_Y));
    OR4 OR4_1408 (.A(OR4_2255_Y), .B(OR4_280_Y), .C(OR4_1994_Y), .D(
        OR4_376_Y), .Y(OR4_1408_Y));
    OR4 OR4_1025 (.A(\A_DOUT_TEMPR16[31] ), .B(\A_DOUT_TEMPR17[31] ), 
        .C(\A_DOUT_TEMPR18[31] ), .D(\A_DOUT_TEMPR19[31] ), .Y(
        OR4_1025_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%82%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R82C5 (
        .A_DOUT({nc8550, nc8551, nc8552, nc8553, nc8554, nc8555, 
        nc8556, nc8557, nc8558, nc8559, nc8560, nc8561, nc8562, nc8563, 
        nc8564, \A_DOUT_TEMPR82[29] , \A_DOUT_TEMPR82[28] , 
        \A_DOUT_TEMPR82[27] , \A_DOUT_TEMPR82[26] , 
        \A_DOUT_TEMPR82[25] }), .B_DOUT({nc8565, nc8566, nc8567, 
        nc8568, nc8569, nc8570, nc8571, nc8572, nc8573, nc8574, nc8575, 
        nc8576, nc8577, nc8578, nc8579, \B_DOUT_TEMPR82[29] , 
        \B_DOUT_TEMPR82[28] , \B_DOUT_TEMPR82[27] , 
        \B_DOUT_TEMPR82[26] , \B_DOUT_TEMPR82[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[82][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_606 (.A(\B_DOUT_TEMPR40[21] ), .B(\B_DOUT_TEMPR41[21] ), 
        .C(\B_DOUT_TEMPR42[21] ), .D(\B_DOUT_TEMPR43[21] ), .Y(
        OR4_606_Y));
    OR4 OR4_2824 (.A(OR4_2947_Y), .B(OR4_2232_Y), .C(OR4_1149_Y), .D(
        OR4_2720_Y), .Y(OR4_2824_Y));
    OR4 OR4_459 (.A(\B_DOUT_TEMPR32[12] ), .B(\B_DOUT_TEMPR33[12] ), 
        .C(\B_DOUT_TEMPR34[12] ), .D(\B_DOUT_TEMPR35[12] ), .Y(
        OR4_459_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%65%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R65C0 (
        .A_DOUT({nc8580, nc8581, nc8582, nc8583, nc8584, nc8585, 
        nc8586, nc8587, nc8588, nc8589, nc8590, nc8591, nc8592, nc8593, 
        nc8594, \A_DOUT_TEMPR65[4] , \A_DOUT_TEMPR65[3] , 
        \A_DOUT_TEMPR65[2] , \A_DOUT_TEMPR65[1] , \A_DOUT_TEMPR65[0] })
        , .B_DOUT({nc8595, nc8596, nc8597, nc8598, nc8599, nc8600, 
        nc8601, nc8602, nc8603, nc8604, nc8605, nc8606, nc8607, nc8608, 
        nc8609, \B_DOUT_TEMPR65[4] , \B_DOUT_TEMPR65[3] , 
        \B_DOUT_TEMPR65[2] , \B_DOUT_TEMPR65[1] , \B_DOUT_TEMPR65[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[65][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[16] , \BLKX1[0] , A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_318 (.A(\B_DOUT_TEMPR91[19] ), .B(\B_DOUT_TEMPR92[19] ), 
        .C(\B_DOUT_TEMPR93[19] ), .D(\B_DOUT_TEMPR94[19] ), .Y(
        OR4_318_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%55%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R55C7 (
        .A_DOUT({nc8610, nc8611, nc8612, nc8613, nc8614, nc8615, 
        nc8616, nc8617, nc8618, nc8619, nc8620, nc8621, nc8622, nc8623, 
        nc8624, \A_DOUT_TEMPR55[39] , \A_DOUT_TEMPR55[38] , 
        \A_DOUT_TEMPR55[37] , \A_DOUT_TEMPR55[36] , 
        \A_DOUT_TEMPR55[35] }), .B_DOUT({nc8625, nc8626, nc8627, 
        nc8628, nc8629, nc8630, nc8631, nc8632, nc8633, nc8634, nc8635, 
        nc8636, nc8637, nc8638, nc8639, \B_DOUT_TEMPR55[39] , 
        \B_DOUT_TEMPR55[38] , \B_DOUT_TEMPR55[37] , 
        \B_DOUT_TEMPR55[36] , \B_DOUT_TEMPR55[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[55][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1299 (.A(\A_DOUT_TEMPR20[6] ), .B(\A_DOUT_TEMPR21[6] ), .C(
        \A_DOUT_TEMPR22[6] ), .D(\A_DOUT_TEMPR23[6] ), .Y(OR4_1299_Y));
    OR4 OR4_3022 (.A(\B_DOUT_TEMPR95[35] ), .B(\B_DOUT_TEMPR96[35] ), 
        .C(\B_DOUT_TEMPR97[35] ), .D(\B_DOUT_TEMPR98[35] ), .Y(
        OR4_3022_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%82%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R82C1 (
        .A_DOUT({nc8640, nc8641, nc8642, nc8643, nc8644, nc8645, 
        nc8646, nc8647, nc8648, nc8649, nc8650, nc8651, nc8652, nc8653, 
        nc8654, \A_DOUT_TEMPR82[9] , \A_DOUT_TEMPR82[8] , 
        \A_DOUT_TEMPR82[7] , \A_DOUT_TEMPR82[6] , \A_DOUT_TEMPR82[5] })
        , .B_DOUT({nc8655, nc8656, nc8657, nc8658, nc8659, nc8660, 
        nc8661, nc8662, nc8663, nc8664, nc8665, nc8666, nc8667, nc8668, 
        nc8669, \B_DOUT_TEMPR82[9] , \B_DOUT_TEMPR82[8] , 
        \B_DOUT_TEMPR82[7] , \B_DOUT_TEMPR82[6] , \B_DOUT_TEMPR82[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[82][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_426 (.A(\A_DOUT_TEMPR8[31] ), .B(\A_DOUT_TEMPR9[31] ), .C(
        \A_DOUT_TEMPR10[31] ), .D(\A_DOUT_TEMPR11[31] ), .Y(OR4_426_Y));
    OR4 OR4_715 (.A(OR4_1743_Y), .B(OR4_693_Y), .C(OR4_2336_Y), .D(
        OR4_287_Y), .Y(OR4_715_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%102%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R102C1 (
        .A_DOUT({nc8670, nc8671, nc8672, nc8673, nc8674, nc8675, 
        nc8676, nc8677, nc8678, nc8679, nc8680, nc8681, nc8682, nc8683, 
        nc8684, \A_DOUT_TEMPR102[9] , \A_DOUT_TEMPR102[8] , 
        \A_DOUT_TEMPR102[7] , \A_DOUT_TEMPR102[6] , 
        \A_DOUT_TEMPR102[5] }), .B_DOUT({nc8685, nc8686, nc8687, 
        nc8688, nc8689, nc8690, nc8691, nc8692, nc8693, nc8694, nc8695, 
        nc8696, nc8697, nc8698, nc8699, \B_DOUT_TEMPR102[9] , 
        \B_DOUT_TEMPR102[8] , \B_DOUT_TEMPR102[7] , 
        \B_DOUT_TEMPR102[6] , \B_DOUT_TEMPR102[5] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[102][1] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[9], 
        B_DIN[8], B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1169 (.A(\A_DOUT_TEMPR64[14] ), .B(\A_DOUT_TEMPR65[14] ), 
        .C(\A_DOUT_TEMPR66[14] ), .D(\A_DOUT_TEMPR67[14] ), .Y(
        OR4_1169_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%24%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R24C7 (
        .A_DOUT({nc8700, nc8701, nc8702, nc8703, nc8704, nc8705, 
        nc8706, nc8707, nc8708, nc8709, nc8710, nc8711, nc8712, nc8713, 
        nc8714, \A_DOUT_TEMPR24[39] , \A_DOUT_TEMPR24[38] , 
        \A_DOUT_TEMPR24[37] , \A_DOUT_TEMPR24[36] , 
        \A_DOUT_TEMPR24[35] }), .B_DOUT({nc8715, nc8716, nc8717, 
        nc8718, nc8719, nc8720, nc8721, nc8722, nc8723, nc8724, nc8725, 
        nc8726, nc8727, nc8728, nc8729, \B_DOUT_TEMPR24[39] , 
        \B_DOUT_TEMPR24[38] , \B_DOUT_TEMPR24[37] , 
        \B_DOUT_TEMPR24[36] , \B_DOUT_TEMPR24[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[24][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2944 (.A(\A_DOUT_TEMPR64[26] ), .B(\A_DOUT_TEMPR65[26] ), 
        .C(\A_DOUT_TEMPR66[26] ), .D(\A_DOUT_TEMPR67[26] ), .Y(
        OR4_2944_Y));
    OR4 OR4_2034 (.A(\A_DOUT_TEMPR4[16] ), .B(\A_DOUT_TEMPR5[16] ), .C(
        \A_DOUT_TEMPR6[16] ), .D(\A_DOUT_TEMPR7[16] ), .Y(OR4_2034_Y));
    OR4 OR4_1500 (.A(OR4_954_Y), .B(OR4_1245_Y), .C(OR4_879_Y), .D(
        OR4_1261_Y), .Y(OR4_1500_Y));
    OR4 OR4_2036 (.A(\B_DOUT_TEMPR32[35] ), .B(\B_DOUT_TEMPR33[35] ), 
        .C(\B_DOUT_TEMPR34[35] ), .D(\B_DOUT_TEMPR35[35] ), .Y(
        OR4_2036_Y));
    OR4 OR4_1827 (.A(\A_DOUT_TEMPR32[3] ), .B(\A_DOUT_TEMPR33[3] ), .C(
        \A_DOUT_TEMPR34[3] ), .D(\A_DOUT_TEMPR35[3] ), .Y(OR4_1827_Y));
    OR4 OR4_3014 (.A(\A_DOUT_TEMPR44[37] ), .B(\A_DOUT_TEMPR45[37] ), 
        .C(\A_DOUT_TEMPR46[37] ), .D(\A_DOUT_TEMPR47[37] ), .Y(
        OR4_3014_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%37%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R37C5 (
        .A_DOUT({nc8730, nc8731, nc8732, nc8733, nc8734, nc8735, 
        nc8736, nc8737, nc8738, nc8739, nc8740, nc8741, nc8742, nc8743, 
        nc8744, \A_DOUT_TEMPR37[29] , \A_DOUT_TEMPR37[28] , 
        \A_DOUT_TEMPR37[27] , \A_DOUT_TEMPR37[26] , 
        \A_DOUT_TEMPR37[25] }), .B_DOUT({nc8745, nc8746, nc8747, 
        nc8748, nc8749, nc8750, nc8751, nc8752, nc8753, nc8754, nc8755, 
        nc8756, nc8757, nc8758, nc8759, \B_DOUT_TEMPR37[29] , 
        \B_DOUT_TEMPR37[28] , \B_DOUT_TEMPR37[27] , 
        \B_DOUT_TEMPR37[26] , \B_DOUT_TEMPR37[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[37][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_939 (.A(\A_DOUT_TEMPR24[3] ), .B(\A_DOUT_TEMPR25[3] ), .C(
        \A_DOUT_TEMPR26[3] ), .D(\A_DOUT_TEMPR27[3] ), .Y(OR4_939_Y));
    OR4 OR4_3016 (.A(\A_DOUT_TEMPR20[13] ), .B(\A_DOUT_TEMPR21[13] ), 
        .C(\A_DOUT_TEMPR22[13] ), .D(\A_DOUT_TEMPR23[13] ), .Y(
        OR4_3016_Y));
    OR4 OR4_1034 (.A(\A_DOUT_TEMPR32[26] ), .B(\A_DOUT_TEMPR33[26] ), 
        .C(\A_DOUT_TEMPR34[26] ), .D(\A_DOUT_TEMPR35[26] ), .Y(
        OR4_1034_Y));
    OR4 OR4_2908 (.A(\A_DOUT_TEMPR32[11] ), .B(\A_DOUT_TEMPR33[11] ), 
        .C(\A_DOUT_TEMPR34[11] ), .D(\A_DOUT_TEMPR35[11] ), .Y(
        OR4_2908_Y));
    OR4 OR4_2946 (.A(OR4_678_Y), .B(OR4_1650_Y), .C(OR4_2332_Y), .D(
        OR4_995_Y), .Y(OR4_2946_Y));
    OR4 OR4_1036 (.A(OR4_1208_Y), .B(OR4_2891_Y), .C(OR4_2292_Y), .D(
        OR4_590_Y), .Y(OR4_1036_Y));
    OR4 OR4_2576 (.A(OR4_399_Y), .B(OR4_2636_Y), .C(OR4_1596_Y), .D(
        OR4_1902_Y), .Y(OR4_2576_Y));
    OR4 OR4_2564 (.A(\A_DOUT_TEMPR75[20] ), .B(\A_DOUT_TEMPR76[20] ), 
        .C(\A_DOUT_TEMPR77[20] ), .D(\A_DOUT_TEMPR78[20] ), .Y(
        OR4_2564_Y));
    OR4 OR4_2777 (.A(\A_DOUT_TEMPR91[3] ), .B(\A_DOUT_TEMPR92[3] ), .C(
        \A_DOUT_TEMPR93[3] ), .D(\A_DOUT_TEMPR94[3] ), .Y(OR4_2777_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%73%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R73C0 (
        .A_DOUT({nc8760, nc8761, nc8762, nc8763, nc8764, nc8765, 
        nc8766, nc8767, nc8768, nc8769, nc8770, nc8771, nc8772, nc8773, 
        nc8774, \A_DOUT_TEMPR73[4] , \A_DOUT_TEMPR73[3] , 
        \A_DOUT_TEMPR73[2] , \A_DOUT_TEMPR73[1] , \A_DOUT_TEMPR73[0] })
        , .B_DOUT({nc8775, nc8776, nc8777, nc8778, nc8779, nc8780, 
        nc8781, nc8782, nc8783, nc8784, nc8785, nc8786, nc8787, nc8788, 
        nc8789, \B_DOUT_TEMPR73[4] , \B_DOUT_TEMPR73[3] , 
        \B_DOUT_TEMPR73[2] , \B_DOUT_TEMPR73[1] , \B_DOUT_TEMPR73[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[73][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_151 (.A(\B_DOUT_TEMPR0[16] ), .B(\B_DOUT_TEMPR1[16] ), .C(
        \B_DOUT_TEMPR2[16] ), .D(\B_DOUT_TEMPR3[16] ), .Y(OR4_151_Y));
    OR4 OR4_2571 (.A(OR4_1042_Y), .B(OR4_2595_Y), .C(OR4_370_Y), .D(
        OR4_2425_Y), .Y(OR4_2571_Y));
    OR4 OR4_104 (.A(\A_DOUT_TEMPR16[37] ), .B(\A_DOUT_TEMPR17[37] ), 
        .C(\A_DOUT_TEMPR18[37] ), .D(\A_DOUT_TEMPR19[37] ), .Y(
        OR4_104_Y));
    OR4 OR4_304 (.A(\A_DOUT_TEMPR60[39] ), .B(\A_DOUT_TEMPR61[39] ), 
        .C(\A_DOUT_TEMPR62[39] ), .D(\A_DOUT_TEMPR63[39] ), .Y(
        OR4_304_Y));
    OR4 OR4_2333 (.A(OR4_598_Y), .B(OR4_917_Y), .C(OR4_535_Y), .D(
        OR4_947_Y), .Y(OR4_2333_Y));
    OR4 OR4_918 (.A(\A_DOUT_TEMPR68[3] ), .B(\A_DOUT_TEMPR69[3] ), .C(
        \A_DOUT_TEMPR70[3] ), .D(\A_DOUT_TEMPR71[3] ), .Y(OR4_918_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%103%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R103C1 (
        .A_DOUT({nc8790, nc8791, nc8792, nc8793, nc8794, nc8795, 
        nc8796, nc8797, nc8798, nc8799, nc8800, nc8801, nc8802, nc8803, 
        nc8804, \A_DOUT_TEMPR103[9] , \A_DOUT_TEMPR103[8] , 
        \A_DOUT_TEMPR103[7] , \A_DOUT_TEMPR103[6] , 
        \A_DOUT_TEMPR103[5] }), .B_DOUT({nc8805, nc8806, nc8807, 
        nc8808, nc8809, nc8810, nc8811, nc8812, nc8813, nc8814, nc8815, 
        nc8816, nc8817, nc8818, nc8819, \B_DOUT_TEMPR103[9] , 
        \B_DOUT_TEMPR103[8] , \B_DOUT_TEMPR103[7] , 
        \B_DOUT_TEMPR103[6] , \B_DOUT_TEMPR103[5] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[103][1] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[9], 
        B_DIN[8], B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_33 (.A(\A_DOUT_TEMPR36[29] ), .B(\A_DOUT_TEMPR37[29] ), .C(
        \A_DOUT_TEMPR38[29] ), .D(\A_DOUT_TEMPR39[29] ), .Y(OR4_33_Y));
    OR4 OR4_1333 (.A(OR4_555_Y), .B(OR4_963_Y), .C(OR4_1672_Y), .D(
        OR4_2496_Y), .Y(OR4_1333_Y));
    OR4 OR4_1556 (.A(\B_DOUT_TEMPR48[11] ), .B(\B_DOUT_TEMPR49[11] ), 
        .C(\B_DOUT_TEMPR50[11] ), .D(\B_DOUT_TEMPR51[11] ), .Y(
        OR4_1556_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKY1[0]  (.A(B_ADDR[13]), .Y(
        \BLKY1[0] ));
    OR4 OR4_1757 (.A(OR4_90_Y), .B(OR4_1300_Y), .C(OR4_2320_Y), .D(
        OR4_993_Y), .Y(OR4_1757_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%77%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R77C7 (
        .A_DOUT({nc8820, nc8821, nc8822, nc8823, nc8824, nc8825, 
        nc8826, nc8827, nc8828, nc8829, nc8830, nc8831, nc8832, nc8833, 
        nc8834, \A_DOUT_TEMPR77[39] , \A_DOUT_TEMPR77[38] , 
        \A_DOUT_TEMPR77[37] , \A_DOUT_TEMPR77[36] , 
        \A_DOUT_TEMPR77[35] }), .B_DOUT({nc8835, nc8836, nc8837, 
        nc8838, nc8839, nc8840, nc8841, nc8842, nc8843, nc8844, nc8845, 
        nc8846, nc8847, nc8848, nc8849, \B_DOUT_TEMPR77[39] , 
        \B_DOUT_TEMPR77[38] , \B_DOUT_TEMPR77[37] , 
        \B_DOUT_TEMPR77[36] , \B_DOUT_TEMPR77[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[77][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR2 OR2_79 (.A(\B_DOUT_TEMPR72[20] ), .B(\B_DOUT_TEMPR73[20] ), .Y(
        OR2_79_Y));
    OR4 OR4_1385 (.A(\B_DOUT_TEMPR32[3] ), .B(\B_DOUT_TEMPR33[3] ), .C(
        \B_DOUT_TEMPR34[3] ), .D(\B_DOUT_TEMPR35[3] ), .Y(OR4_1385_Y));
    OR4 OR4_1551 (.A(\B_DOUT_TEMPR0[17] ), .B(\B_DOUT_TEMPR1[17] ), .C(
        \B_DOUT_TEMPR2[17] ), .D(\B_DOUT_TEMPR3[17] ), .Y(OR4_1551_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%69%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R69C1 (
        .A_DOUT({nc8850, nc8851, nc8852, nc8853, nc8854, nc8855, 
        nc8856, nc8857, nc8858, nc8859, nc8860, nc8861, nc8862, nc8863, 
        nc8864, \A_DOUT_TEMPR69[9] , \A_DOUT_TEMPR69[8] , 
        \A_DOUT_TEMPR69[7] , \A_DOUT_TEMPR69[6] , \A_DOUT_TEMPR69[5] })
        , .B_DOUT({nc8865, nc8866, nc8867, nc8868, nc8869, nc8870, 
        nc8871, nc8872, nc8873, nc8874, nc8875, nc8876, nc8877, nc8878, 
        nc8879, \B_DOUT_TEMPR69[9] , \B_DOUT_TEMPR69[8] , 
        \B_DOUT_TEMPR69[7] , \B_DOUT_TEMPR69[6] , \B_DOUT_TEMPR69[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[69][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_876 (.A(\B_DOUT_TEMPR60[22] ), .B(\B_DOUT_TEMPR61[22] ), 
        .C(\B_DOUT_TEMPR62[22] ), .D(\B_DOUT_TEMPR63[22] ), .Y(
        OR4_876_Y));
    OR4 OR4_1905 (.A(\B_DOUT_TEMPR64[9] ), .B(\B_DOUT_TEMPR65[9] ), .C(
        \B_DOUT_TEMPR66[9] ), .D(\B_DOUT_TEMPR67[9] ), .Y(OR4_1905_Y));
    OR4 OR4_118 (.A(\A_DOUT_TEMPR48[13] ), .B(\A_DOUT_TEMPR49[13] ), 
        .C(\A_DOUT_TEMPR50[13] ), .D(\A_DOUT_TEMPR51[13] ), .Y(
        OR4_118_Y));
    OR4 OR4_2261 (.A(OR4_1606_Y), .B(OR4_328_Y), .C(OR4_1055_Y), .D(
        OR4_1349_Y), .Y(OR4_2261_Y));
    OR4 OR4_2107 (.A(\A_DOUT_TEMPR32[23] ), .B(\A_DOUT_TEMPR33[23] ), 
        .C(\A_DOUT_TEMPR34[23] ), .D(\A_DOUT_TEMPR35[23] ), .Y(
        OR4_2107_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%35%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R35C7 (
        .A_DOUT({nc8880, nc8881, nc8882, nc8883, nc8884, nc8885, 
        nc8886, nc8887, nc8888, nc8889, nc8890, nc8891, nc8892, nc8893, 
        nc8894, \A_DOUT_TEMPR35[39] , \A_DOUT_TEMPR35[38] , 
        \A_DOUT_TEMPR35[37] , \A_DOUT_TEMPR35[36] , 
        \A_DOUT_TEMPR35[35] }), .B_DOUT({nc8895, nc8896, nc8897, 
        nc8898, nc8899, nc8900, nc8901, nc8902, nc8903, nc8904, nc8905, 
        nc8906, nc8907, nc8908, nc8909, \B_DOUT_TEMPR35[39] , 
        \B_DOUT_TEMPR35[38] , \B_DOUT_TEMPR35[37] , 
        \B_DOUT_TEMPR35[36] , \B_DOUT_TEMPR35[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[35][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_255 (.A(OR4_212_Y), .B(OR4_2641_Y), .C(OR4_1093_Y), .D(
        OR4_2642_Y), .Y(OR4_255_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%18%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R18C0 (
        .A_DOUT({nc8910, nc8911, nc8912, nc8913, nc8914, nc8915, 
        nc8916, nc8917, nc8918, nc8919, nc8920, nc8921, nc8922, nc8923, 
        nc8924, \A_DOUT_TEMPR18[4] , \A_DOUT_TEMPR18[3] , 
        \A_DOUT_TEMPR18[2] , \A_DOUT_TEMPR18[1] , \A_DOUT_TEMPR18[0] })
        , .B_DOUT({nc8925, nc8926, nc8927, nc8928, nc8929, nc8930, 
        nc8931, nc8932, nc8933, nc8934, nc8935, nc8936, nc8937, nc8938, 
        nc8939, \B_DOUT_TEMPR18[4] , \B_DOUT_TEMPR18[3] , 
        \B_DOUT_TEMPR18[2] , \B_DOUT_TEMPR18[1] , \B_DOUT_TEMPR18[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[18][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2604 (.A(\A_DOUT_TEMPR75[34] ), .B(\A_DOUT_TEMPR76[34] ), 
        .C(\A_DOUT_TEMPR77[34] ), .D(\A_DOUT_TEMPR78[34] ), .Y(
        OR4_2604_Y));
    OR4 OR4_370 (.A(\A_DOUT_TEMPR8[15] ), .B(\A_DOUT_TEMPR9[15] ), .C(
        \A_DOUT_TEMPR10[15] ), .D(\A_DOUT_TEMPR11[15] ), .Y(OR4_370_Y));
    OR4 OR4_319 (.A(OR4_1781_Y), .B(OR4_3001_Y), .C(OR4_2563_Y), .D(
        OR4_1218_Y), .Y(OR4_319_Y));
    OR4 OR4_1609 (.A(\A_DOUT_TEMPR60[15] ), .B(\A_DOUT_TEMPR61[15] ), 
        .C(\A_DOUT_TEMPR62[15] ), .D(\A_DOUT_TEMPR63[15] ), .Y(
        OR4_1609_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%69%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R69C2 (
        .A_DOUT({nc8940, nc8941, nc8942, nc8943, nc8944, nc8945, 
        nc8946, nc8947, nc8948, nc8949, nc8950, nc8951, nc8952, nc8953, 
        nc8954, \A_DOUT_TEMPR69[14] , \A_DOUT_TEMPR69[13] , 
        \A_DOUT_TEMPR69[12] , \A_DOUT_TEMPR69[11] , 
        \A_DOUT_TEMPR69[10] }), .B_DOUT({nc8955, nc8956, nc8957, 
        nc8958, nc8959, nc8960, nc8961, nc8962, nc8963, nc8964, nc8965, 
        nc8966, nc8967, nc8968, nc8969, \B_DOUT_TEMPR69[14] , 
        \B_DOUT_TEMPR69[13] , \B_DOUT_TEMPR69[12] , 
        \B_DOUT_TEMPR69[11] , \B_DOUT_TEMPR69[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[69][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_446 (.A(OR4_1920_Y), .B(OR4_35_Y), .C(OR4_384_Y), .D(
        OR4_828_Y), .Y(OR4_446_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%65%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R65C1 (
        .A_DOUT({nc8970, nc8971, nc8972, nc8973, nc8974, nc8975, 
        nc8976, nc8977, nc8978, nc8979, nc8980, nc8981, nc8982, nc8983, 
        nc8984, \A_DOUT_TEMPR65[9] , \A_DOUT_TEMPR65[8] , 
        \A_DOUT_TEMPR65[7] , \A_DOUT_TEMPR65[6] , \A_DOUT_TEMPR65[5] })
        , .B_DOUT({nc8985, nc8986, nc8987, nc8988, nc8989, nc8990, 
        nc8991, nc8992, nc8993, nc8994, nc8995, nc8996, nc8997, nc8998, 
        nc8999, \B_DOUT_TEMPR65[9] , \B_DOUT_TEMPR65[8] , 
        \B_DOUT_TEMPR65[7] , \B_DOUT_TEMPR65[6] , \B_DOUT_TEMPR65[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[65][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[16] , \BLKX1[0] , A_ADDR[12]}), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], 
        A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%116%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R116C1 (
        .A_DOUT({nc9000, nc9001, nc9002, nc9003, nc9004, nc9005, 
        nc9006, nc9007, nc9008, nc9009, nc9010, nc9011, nc9012, nc9013, 
        nc9014, \A_DOUT_TEMPR116[9] , \A_DOUT_TEMPR116[8] , 
        \A_DOUT_TEMPR116[7] , \A_DOUT_TEMPR116[6] , 
        \A_DOUT_TEMPR116[5] }), .B_DOUT({nc9015, nc9016, nc9017, 
        nc9018, nc9019, nc9020, nc9021, nc9022, nc9023, nc9024, nc9025, 
        nc9026, nc9027, nc9028, nc9029, \B_DOUT_TEMPR116[9] , 
        \B_DOUT_TEMPR116[8] , \B_DOUT_TEMPR116[7] , 
        \B_DOUT_TEMPR116[6] , \B_DOUT_TEMPR116[5] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[116][1] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(
        A_REN), .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[9], 
        B_DIN[8], B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({
        GND, \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%57%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R57C2 (
        .A_DOUT({nc9030, nc9031, nc9032, nc9033, nc9034, nc9035, 
        nc9036, nc9037, nc9038, nc9039, nc9040, nc9041, nc9042, nc9043, 
        nc9044, \A_DOUT_TEMPR57[14] , \A_DOUT_TEMPR57[13] , 
        \A_DOUT_TEMPR57[12] , \A_DOUT_TEMPR57[11] , 
        \A_DOUT_TEMPR57[10] }), .B_DOUT({nc9045, nc9046, nc9047, 
        nc9048, nc9049, nc9050, nc9051, nc9052, nc9053, nc9054, nc9055, 
        nc9056, nc9057, nc9058, nc9059, \B_DOUT_TEMPR57[14] , 
        \B_DOUT_TEMPR57[13] , \B_DOUT_TEMPR57[12] , 
        \B_DOUT_TEMPR57[11] , \B_DOUT_TEMPR57[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[57][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_656 (.A(\A_DOUT_TEMPR0[36] ), .B(\A_DOUT_TEMPR1[36] ), .C(
        \A_DOUT_TEMPR2[36] ), .D(\A_DOUT_TEMPR3[36] ), .Y(OR4_656_Y));
    OR2 OR2_42 (.A(\A_DOUT_TEMPR72[20] ), .B(\A_DOUT_TEMPR73[20] ), .Y(
        OR2_42_Y));
    OR4 OR4_2615 (.A(\A_DOUT_TEMPR44[0] ), .B(\A_DOUT_TEMPR45[0] ), .C(
        \A_DOUT_TEMPR46[0] ), .D(\A_DOUT_TEMPR47[0] ), .Y(OR4_2615_Y));
    OR4 OR4_1862 (.A(\A_DOUT_TEMPR48[26] ), .B(\A_DOUT_TEMPR49[26] ), 
        .C(\A_DOUT_TEMPR50[26] ), .D(\A_DOUT_TEMPR51[26] ), .Y(
        OR4_1862_Y));
    OR4 OR4_2325 (.A(OR4_691_Y), .B(OR4_1344_Y), .C(OR4_912_Y), .D(
        OR4_2582_Y), .Y(OR4_2325_Y));
    OR4 OR4_499 (.A(\B_DOUT_TEMPR4[7] ), .B(\B_DOUT_TEMPR5[7] ), .C(
        \B_DOUT_TEMPR6[7] ), .D(\B_DOUT_TEMPR7[7] ), .Y(OR4_499_Y));
    OR4 OR4_212 (.A(OR4_37_Y), .B(OR4_1241_Y), .C(OR2_52_Y), .D(
        \A_DOUT_TEMPR74[13] ), .Y(OR4_212_Y));
    OR4 OR4_806 (.A(\B_DOUT_TEMPR95[26] ), .B(\B_DOUT_TEMPR96[26] ), 
        .C(\B_DOUT_TEMPR97[26] ), .D(\B_DOUT_TEMPR98[26] ), .Y(
        OR4_806_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%94%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R94C0 (
        .A_DOUT({nc9060, nc9061, nc9062, nc9063, nc9064, nc9065, 
        nc9066, nc9067, nc9068, nc9069, nc9070, nc9071, nc9072, nc9073, 
        nc9074, \A_DOUT_TEMPR94[4] , \A_DOUT_TEMPR94[3] , 
        \A_DOUT_TEMPR94[2] , \A_DOUT_TEMPR94[1] , \A_DOUT_TEMPR94[0] })
        , .B_DOUT({nc9075, nc9076, nc9077, nc9078, nc9079, nc9080, 
        nc9081, nc9082, nc9083, nc9084, nc9085, nc9086, nc9087, nc9088, 
        nc9089, \B_DOUT_TEMPR94[4] , \B_DOUT_TEMPR94[3] , 
        \B_DOUT_TEMPR94[2] , \B_DOUT_TEMPR94[1] , \B_DOUT_TEMPR94[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[94][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_83 (.A(OR4_2103_Y), .B(OR4_1584_Y), .C(OR4_40_Y), .D(
        OR4_1585_Y), .Y(OR4_83_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%15%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R15C0 (
        .A_DOUT({nc9090, nc9091, nc9092, nc9093, nc9094, nc9095, 
        nc9096, nc9097, nc9098, nc9099, nc9100, nc9101, nc9102, nc9103, 
        nc9104, \A_DOUT_TEMPR15[4] , \A_DOUT_TEMPR15[3] , 
        \A_DOUT_TEMPR15[2] , \A_DOUT_TEMPR15[1] , \A_DOUT_TEMPR15[0] })
        , .B_DOUT({nc9105, nc9106, nc9107, nc9108, nc9109, nc9110, 
        nc9111, nc9112, nc9113, nc9114, nc9115, nc9116, nc9117, nc9118, 
        nc9119, \B_DOUT_TEMPR15[4] , \B_DOUT_TEMPR15[3] , 
        \B_DOUT_TEMPR15[2] , \B_DOUT_TEMPR15[1] , \B_DOUT_TEMPR15[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[15][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[3] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], 
        A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_300 (.A(\A_DOUT_TEMPR79[3] ), .B(\A_DOUT_TEMPR80[3] ), .C(
        \A_DOUT_TEMPR81[3] ), .D(\A_DOUT_TEMPR82[3] ), .Y(OR4_300_Y));
    OR4 OR4_368 (.A(OR4_2208_Y), .B(OR4_2041_Y), .C(OR4_2935_Y), .D(
        OR4_1086_Y), .Y(OR4_368_Y));
    OR4 OR4_2617 (.A(\B_DOUT_TEMPR52[13] ), .B(\B_DOUT_TEMPR53[13] ), 
        .C(\B_DOUT_TEMPR54[13] ), .D(\B_DOUT_TEMPR55[13] ), .Y(
        OR4_2617_Y));
    OR4 OR4_154 (.A(\A_DOUT_TEMPR28[34] ), .B(\A_DOUT_TEMPR29[34] ), 
        .C(\A_DOUT_TEMPR30[34] ), .D(\A_DOUT_TEMPR31[34] ), .Y(
        OR4_154_Y));
    OR4 OR4_354 (.A(\B_DOUT_TEMPR79[15] ), .B(\B_DOUT_TEMPR80[15] ), 
        .C(\B_DOUT_TEMPR81[15] ), .D(\B_DOUT_TEMPR82[15] ), .Y(
        OR4_354_Y));
    OR4 OR4_765 (.A(\A_DOUT_TEMPR36[19] ), .B(\A_DOUT_TEMPR37[19] ), 
        .C(\A_DOUT_TEMPR38[19] ), .D(\A_DOUT_TEMPR39[19] ), .Y(
        OR4_765_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%23%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R23C4 (
        .A_DOUT({nc9120, nc9121, nc9122, nc9123, nc9124, nc9125, 
        nc9126, nc9127, nc9128, nc9129, nc9130, nc9131, nc9132, nc9133, 
        nc9134, \A_DOUT_TEMPR23[24] , \A_DOUT_TEMPR23[23] , 
        \A_DOUT_TEMPR23[22] , \A_DOUT_TEMPR23[21] , 
        \A_DOUT_TEMPR23[20] }), .B_DOUT({nc9135, nc9136, nc9137, 
        nc9138, nc9139, nc9140, nc9141, nc9142, nc9143, nc9144, nc9145, 
        nc9146, nc9147, nc9148, nc9149, \B_DOUT_TEMPR23[24] , 
        \B_DOUT_TEMPR23[23] , \B_DOUT_TEMPR23[22] , 
        \B_DOUT_TEMPR23[21] , \B_DOUT_TEMPR23[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[23][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1663 (.A(\B_DOUT_TEMPR44[33] ), .B(\B_DOUT_TEMPR45[33] ), 
        .C(\B_DOUT_TEMPR46[33] ), .D(\B_DOUT_TEMPR47[33] ), .Y(
        OR4_1663_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_0 (.A(A_ADDR[16]), .B(A_ADDR[15]), .C(
        A_ADDR[14]), .Y(CFG3_0_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%96%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R96C7 (
        .A_DOUT({nc9150, nc9151, nc9152, nc9153, nc9154, nc9155, 
        nc9156, nc9157, nc9158, nc9159, nc9160, nc9161, nc9162, nc9163, 
        nc9164, \A_DOUT_TEMPR96[39] , \A_DOUT_TEMPR96[38] , 
        \A_DOUT_TEMPR96[37] , \A_DOUT_TEMPR96[36] , 
        \A_DOUT_TEMPR96[35] }), .B_DOUT({nc9165, nc9166, nc9167, 
        nc9168, nc9169, nc9170, nc9171, nc9172, nc9173, nc9174, nc9175, 
        nc9176, nc9177, nc9178, nc9179, \B_DOUT_TEMPR96[39] , 
        \B_DOUT_TEMPR96[38] , \B_DOUT_TEMPR96[37] , 
        \B_DOUT_TEMPR96[36] , \B_DOUT_TEMPR96[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[96][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%67%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R67C5 (
        .A_DOUT({nc9180, nc9181, nc9182, nc9183, nc9184, nc9185, 
        nc9186, nc9187, nc9188, nc9189, nc9190, nc9191, nc9192, nc9193, 
        nc9194, \A_DOUT_TEMPR67[29] , \A_DOUT_TEMPR67[28] , 
        \A_DOUT_TEMPR67[27] , \A_DOUT_TEMPR67[26] , 
        \A_DOUT_TEMPR67[25] }), .B_DOUT({nc9195, nc9196, nc9197, 
        nc9198, nc9199, nc9200, nc9201, nc9202, nc9203, nc9204, nc9205, 
        nc9206, nc9207, nc9208, nc9209, \B_DOUT_TEMPR67[29] , 
        \B_DOUT_TEMPR67[28] , \B_DOUT_TEMPR67[27] , 
        \B_DOUT_TEMPR67[26] , \B_DOUT_TEMPR67[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[67][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_191 (.A(\B_DOUT_TEMPR64[12] ), .B(\B_DOUT_TEMPR65[12] ), 
        .C(\B_DOUT_TEMPR66[12] ), .D(\B_DOUT_TEMPR67[12] ), .Y(
        OR4_191_Y));
    OR4 OR4_1210 (.A(\A_DOUT_TEMPR111[0] ), .B(\A_DOUT_TEMPR112[0] ), 
        .C(\A_DOUT_TEMPR113[0] ), .D(\A_DOUT_TEMPR114[0] ), .Y(
        OR4_1210_Y));
    OR4 OR4_1969 (.A(\B_DOUT_TEMPR44[6] ), .B(\B_DOUT_TEMPR45[6] ), .C(
        \B_DOUT_TEMPR46[6] ), .D(\B_DOUT_TEMPR47[6] ), .Y(OR4_1969_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%97%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R97C6 (
        .A_DOUT({nc9210, nc9211, nc9212, nc9213, nc9214, nc9215, 
        nc9216, nc9217, nc9218, nc9219, nc9220, nc9221, nc9222, nc9223, 
        nc9224, \A_DOUT_TEMPR97[34] , \A_DOUT_TEMPR97[33] , 
        \A_DOUT_TEMPR97[32] , \A_DOUT_TEMPR97[31] , 
        \A_DOUT_TEMPR97[30] }), .B_DOUT({nc9225, nc9226, nc9227, 
        nc9228, nc9229, nc9230, nc9231, nc9232, nc9233, nc9234, nc9235, 
        nc9236, nc9237, nc9238, nc9239, \B_DOUT_TEMPR97[34] , 
        \B_DOUT_TEMPR97[33] , \B_DOUT_TEMPR97[32] , 
        \B_DOUT_TEMPR97[31] , \B_DOUT_TEMPR97[30] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[97][6] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[34], A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[34], 
        B_DIN[33], B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%37%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R37C2 (
        .A_DOUT({nc9240, nc9241, nc9242, nc9243, nc9244, nc9245, 
        nc9246, nc9247, nc9248, nc9249, nc9250, nc9251, nc9252, nc9253, 
        nc9254, \A_DOUT_TEMPR37[14] , \A_DOUT_TEMPR37[13] , 
        \A_DOUT_TEMPR37[12] , \A_DOUT_TEMPR37[11] , 
        \A_DOUT_TEMPR37[10] }), .B_DOUT({nc9255, nc9256, nc9257, 
        nc9258, nc9259, nc9260, nc9261, nc9262, nc9263, nc9264, nc9265, 
        nc9266, nc9267, nc9268, nc9269, \B_DOUT_TEMPR37[14] , 
        \B_DOUT_TEMPR37[13] , \B_DOUT_TEMPR37[12] , 
        \B_DOUT_TEMPR37[11] , \B_DOUT_TEMPR37[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[37][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2878 (.A(\B_DOUT_TEMPR68[25] ), .B(\B_DOUT_TEMPR69[25] ), 
        .C(\B_DOUT_TEMPR70[25] ), .D(\B_DOUT_TEMPR71[25] ), .Y(
        OR4_2878_Y));
    OR4 OR4_274 (.A(\A_DOUT_TEMPR83[17] ), .B(\A_DOUT_TEMPR84[17] ), 
        .C(\A_DOUT_TEMPR85[17] ), .D(\A_DOUT_TEMPR86[17] ), .Y(
        OR4_274_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%0%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R0C2 (
        .A_DOUT({nc9270, nc9271, nc9272, nc9273, nc9274, nc9275, 
        nc9276, nc9277, nc9278, nc9279, nc9280, nc9281, nc9282, nc9283, 
        nc9284, \A_DOUT_TEMPR0[14] , \A_DOUT_TEMPR0[13] , 
        \A_DOUT_TEMPR0[12] , \A_DOUT_TEMPR0[11] , \A_DOUT_TEMPR0[10] })
        , .B_DOUT({nc9285, nc9286, nc9287, nc9288, nc9289, nc9290, 
        nc9291, nc9292, nc9293, nc9294, nc9295, nc9296, nc9297, nc9298, 
        nc9299, \B_DOUT_TEMPR0[14] , \B_DOUT_TEMPR0[13] , 
        \B_DOUT_TEMPR0[12] , \B_DOUT_TEMPR0[11] , \B_DOUT_TEMPR0[10] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[0][2] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[14], A_DIN[13], A_DIN[12], 
        A_DIN[11], A_DIN[10]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_44 (.A(\A_DOUT_TEMPR72[32] ), .B(\A_DOUT_TEMPR73[32] ), .Y(
        OR2_44_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%101%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R101C2 (
        .A_DOUT({nc9300, nc9301, nc9302, nc9303, nc9304, nc9305, 
        nc9306, nc9307, nc9308, nc9309, nc9310, nc9311, nc9312, nc9313, 
        nc9314, \A_DOUT_TEMPR101[14] , \A_DOUT_TEMPR101[13] , 
        \A_DOUT_TEMPR101[12] , \A_DOUT_TEMPR101[11] , 
        \A_DOUT_TEMPR101[10] }), .B_DOUT({nc9315, nc9316, nc9317, 
        nc9318, nc9319, nc9320, nc9321, nc9322, nc9323, nc9324, nc9325, 
        nc9326, nc9327, nc9328, nc9329, \B_DOUT_TEMPR101[14] , 
        \B_DOUT_TEMPR101[13] , \B_DOUT_TEMPR101[12] , 
        \B_DOUT_TEMPR101[11] , \B_DOUT_TEMPR101[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[101][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%114%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R114C4 (
        .A_DOUT({nc9330, nc9331, nc9332, nc9333, nc9334, nc9335, 
        nc9336, nc9337, nc9338, nc9339, nc9340, nc9341, nc9342, nc9343, 
        nc9344, \A_DOUT_TEMPR114[24] , \A_DOUT_TEMPR114[23] , 
        \A_DOUT_TEMPR114[22] , \A_DOUT_TEMPR114[21] , 
        \A_DOUT_TEMPR114[20] }), .B_DOUT({nc9345, nc9346, nc9347, 
        nc9348, nc9349, nc9350, nc9351, nc9352, nc9353, nc9354, nc9355, 
        nc9356, nc9357, nc9358, nc9359, \B_DOUT_TEMPR114[24] , 
        \B_DOUT_TEMPR114[23] , \B_DOUT_TEMPR114[22] , 
        \B_DOUT_TEMPR114[21] , \B_DOUT_TEMPR114[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[114][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_770 (.A(\B_DOUT_TEMPR20[21] ), .B(\B_DOUT_TEMPR21[21] ), 
        .C(\B_DOUT_TEMPR22[21] ), .D(\B_DOUT_TEMPR23[21] ), .Y(
        OR4_770_Y));
    OR4 OR4_1007 (.A(\B_DOUT_TEMPR48[25] ), .B(\B_DOUT_TEMPR49[25] ), 
        .C(\B_DOUT_TEMPR50[25] ), .D(\B_DOUT_TEMPR51[25] ), .Y(
        OR4_1007_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%92%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R92C4 (
        .A_DOUT({nc9360, nc9361, nc9362, nc9363, nc9364, nc9365, 
        nc9366, nc9367, nc9368, nc9369, nc9370, nc9371, nc9372, nc9373, 
        nc9374, \A_DOUT_TEMPR92[24] , \A_DOUT_TEMPR92[23] , 
        \A_DOUT_TEMPR92[22] , \A_DOUT_TEMPR92[21] , 
        \A_DOUT_TEMPR92[20] }), .B_DOUT({nc9375, nc9376, nc9377, 
        nc9378, nc9379, nc9380, nc9381, nc9382, nc9383, nc9384, nc9385, 
        nc9386, nc9387, nc9388, nc9389, \B_DOUT_TEMPR92[24] , 
        \B_DOUT_TEMPR92[23] , \B_DOUT_TEMPR92[22] , 
        \B_DOUT_TEMPR92[21] , \B_DOUT_TEMPR92[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[92][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_968 (.A(\A_DOUT_TEMPR8[1] ), .B(\A_DOUT_TEMPR9[1] ), .C(
        \A_DOUT_TEMPR10[1] ), .D(\A_DOUT_TEMPR11[1] ), .Y(OR4_968_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[20]  (.A(CFG3_4_Y), .B(CFG3_3_Y)
        , .Y(\BLKX2[20] ));
    OR4 OR4_1991 (.A(\A_DOUT_TEMPR83[3] ), .B(\A_DOUT_TEMPR84[3] ), .C(
        \A_DOUT_TEMPR85[3] ), .D(\A_DOUT_TEMPR86[3] ), .Y(OR4_1991_Y));
    OR4 OR4_1309 (.A(OR4_970_Y), .B(OR4_1543_Y), .C(OR4_2995_Y), .D(
        OR4_907_Y), .Y(OR4_1309_Y));
    OR4 OR4_1764 (.A(\B_DOUT_TEMPR107[20] ), .B(\B_DOUT_TEMPR108[20] ), 
        .C(\B_DOUT_TEMPR109[20] ), .D(\B_DOUT_TEMPR110[20] ), .Y(
        OR4_1764_Y));
    OR4 OR4_2600 (.A(\A_DOUT_TEMPR8[37] ), .B(\A_DOUT_TEMPR9[37] ), .C(
        \A_DOUT_TEMPR10[37] ), .D(\A_DOUT_TEMPR11[37] ), .Y(OR4_2600_Y)
        );
    OR4 OR4_1316 (.A(\B_DOUT_TEMPR60[25] ), .B(\B_DOUT_TEMPR61[25] ), 
        .C(\B_DOUT_TEMPR62[25] ), .D(\B_DOUT_TEMPR63[25] ), .Y(
        OR4_1316_Y));
    OR4 OR4_1207 (.A(\B_DOUT_TEMPR99[26] ), .B(\B_DOUT_TEMPR100[26] ), 
        .C(\B_DOUT_TEMPR101[26] ), .D(\B_DOUT_TEMPR102[26] ), .Y(
        OR4_1207_Y));
    OR4 OR4_295 (.A(\B_DOUT_TEMPR60[14] ), .B(\B_DOUT_TEMPR61[14] ), 
        .C(\B_DOUT_TEMPR62[14] ), .D(\B_DOUT_TEMPR63[14] ), .Y(
        OR4_295_Y));
    OR4 OR4_2250 (.A(OR4_1326_Y), .B(OR4_2202_Y), .C(OR4_1875_Y), .D(
        OR4_323_Y), .Y(OR4_2250_Y));
    OR4 OR4_1461 (.A(\A_DOUT_TEMPR64[4] ), .B(\A_DOUT_TEMPR65[4] ), .C(
        \A_DOUT_TEMPR66[4] ), .D(\A_DOUT_TEMPR67[4] ), .Y(OR4_1461_Y));
    OR4 OR4_1858 (.A(OR4_302_Y), .B(OR4_120_Y), .C(OR2_1_Y), .D(
        \B_DOUT_TEMPR74[37] ), .Y(OR4_1858_Y));
    OR4 OR4_2008 (.A(\B_DOUT_TEMPR44[25] ), .B(\B_DOUT_TEMPR45[25] ), 
        .C(\B_DOUT_TEMPR46[25] ), .D(\B_DOUT_TEMPR47[25] ), .Y(
        OR4_2008_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%19%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R19C1 (
        .A_DOUT({nc9390, nc9391, nc9392, nc9393, nc9394, nc9395, 
        nc9396, nc9397, nc9398, nc9399, nc9400, nc9401, nc9402, nc9403, 
        nc9404, \A_DOUT_TEMPR19[9] , \A_DOUT_TEMPR19[8] , 
        \A_DOUT_TEMPR19[7] , \A_DOUT_TEMPR19[6] , \A_DOUT_TEMPR19[5] })
        , .B_DOUT({nc9405, nc9406, nc9407, nc9408, nc9409, nc9410, 
        nc9411, nc9412, nc9413, nc9414, nc9415, nc9416, nc9417, nc9418, 
        nc9419, \B_DOUT_TEMPR19[9] , \B_DOUT_TEMPR19[8] , 
        \B_DOUT_TEMPR19[7] , \B_DOUT_TEMPR19[6] , \B_DOUT_TEMPR19[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[19][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], 
        A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1900 (.A(\A_DOUT_TEMPR87[7] ), .B(\A_DOUT_TEMPR88[7] ), .C(
        \A_DOUT_TEMPR89[7] ), .D(\A_DOUT_TEMPR90[7] ), .Y(OR4_1900_Y));
    OR4 OR4_220 (.A(\B_DOUT_TEMPR48[18] ), .B(\B_DOUT_TEMPR49[18] ), 
        .C(\B_DOUT_TEMPR50[18] ), .D(\B_DOUT_TEMPR51[18] ), .Y(
        OR4_220_Y));
    OR4 OR4_168 (.A(OR4_983_Y), .B(OR4_167_Y), .C(OR4_2393_Y), .D(
        OR4_1354_Y), .Y(OR4_168_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%21%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R21C4 (
        .A_DOUT({nc9420, nc9421, nc9422, nc9423, nc9424, nc9425, 
        nc9426, nc9427, nc9428, nc9429, nc9430, nc9431, nc9432, nc9433, 
        nc9434, \A_DOUT_TEMPR21[24] , \A_DOUT_TEMPR21[23] , 
        \A_DOUT_TEMPR21[22] , \A_DOUT_TEMPR21[21] , 
        \A_DOUT_TEMPR21[20] }), .B_DOUT({nc9435, nc9436, nc9437, 
        nc9438, nc9439, nc9440, nc9441, nc9442, nc9443, nc9444, nc9445, 
        nc9446, nc9447, nc9448, nc9449, \B_DOUT_TEMPR21[24] , 
        \B_DOUT_TEMPR21[23] , \B_DOUT_TEMPR21[22] , 
        \B_DOUT_TEMPR21[21] , \B_DOUT_TEMPR21[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[21][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%65%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R65C7 (
        .A_DOUT({nc9450, nc9451, nc9452, nc9453, nc9454, nc9455, 
        nc9456, nc9457, nc9458, nc9459, nc9460, nc9461, nc9462, nc9463, 
        nc9464, \A_DOUT_TEMPR65[39] , \A_DOUT_TEMPR65[38] , 
        \A_DOUT_TEMPR65[37] , \A_DOUT_TEMPR65[36] , 
        \A_DOUT_TEMPR65[35] }), .B_DOUT({nc9465, nc9466, nc9467, 
        nc9468, nc9469, nc9470, nc9471, nc9472, nc9473, nc9474, nc9475, 
        nc9476, nc9477, nc9478, nc9479, \B_DOUT_TEMPR65[39] , 
        \B_DOUT_TEMPR65[38] , \B_DOUT_TEMPR65[37] , 
        \B_DOUT_TEMPR65[36] , \B_DOUT_TEMPR65[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[65][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_696 (.A(OR4_2259_Y), .B(OR4_2795_Y), .C(OR4_1232_Y), .D(
        OR4_2798_Y), .Y(OR4_696_Y));
    OR4 OR4_620 (.A(OR4_129_Y), .B(OR4_2996_Y), .C(OR4_818_Y), .D(
        OR4_2007_Y), .Y(OR4_620_Y));
    OR4 OR4_2314 (.A(\B_DOUT_TEMPR64[27] ), .B(\B_DOUT_TEMPR65[27] ), 
        .C(\B_DOUT_TEMPR66[27] ), .D(\B_DOUT_TEMPR67[27] ), .Y(
        OR4_2314_Y));
    OR4 OR4_369 (.A(\A_DOUT_TEMPR95[22] ), .B(\A_DOUT_TEMPR96[22] ), 
        .C(\A_DOUT_TEMPR97[22] ), .D(\A_DOUT_TEMPR98[22] ), .Y(
        OR4_369_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%19%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R19C2 (
        .A_DOUT({nc9480, nc9481, nc9482, nc9483, nc9484, nc9485, 
        nc9486, nc9487, nc9488, nc9489, nc9490, nc9491, nc9492, nc9493, 
        nc9494, \A_DOUT_TEMPR19[14] , \A_DOUT_TEMPR19[13] , 
        \A_DOUT_TEMPR19[12] , \A_DOUT_TEMPR19[11] , 
        \A_DOUT_TEMPR19[10] }), .B_DOUT({nc9495, nc9496, nc9497, 
        nc9498, nc9499, nc9500, nc9501, nc9502, nc9503, nc9504, nc9505, 
        nc9506, nc9507, nc9508, nc9509, \B_DOUT_TEMPR19[14] , 
        \B_DOUT_TEMPR19[13] , \B_DOUT_TEMPR19[12] , 
        \B_DOUT_TEMPR19[11] , \B_DOUT_TEMPR19[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[19][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[27]  (.A(OR4_2056_Y), .B(OR4_2_Y), .C(OR4_98_Y), 
        .D(OR4_3035_Y), .Y(B_DOUT[27]));
    OR4 OR4_2099 (.A(\B_DOUT_TEMPR0[13] ), .B(\B_DOUT_TEMPR1[13] ), .C(
        \B_DOUT_TEMPR2[13] ), .D(\B_DOUT_TEMPR3[13] ), .Y(OR4_2099_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%15%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R15C1 (
        .A_DOUT({nc9510, nc9511, nc9512, nc9513, nc9514, nc9515, 
        nc9516, nc9517, nc9518, nc9519, nc9520, nc9521, nc9522, nc9523, 
        nc9524, \A_DOUT_TEMPR15[9] , \A_DOUT_TEMPR15[8] , 
        \A_DOUT_TEMPR15[7] , \A_DOUT_TEMPR15[6] , \A_DOUT_TEMPR15[5] })
        , .B_DOUT({nc9525, nc9526, nc9527, nc9528, nc9529, nc9530, 
        nc9531, nc9532, nc9533, nc9534, nc9535, nc9536, nc9537, nc9538, 
        nc9539, \B_DOUT_TEMPR15[9] , \B_DOUT_TEMPR15[8] , 
        \B_DOUT_TEMPR15[7] , \B_DOUT_TEMPR15[6] , \B_DOUT_TEMPR15[5] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[15][1] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[3] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], 
        A_DIN[6], A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%103%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R103C4 (
        .A_DOUT({nc9540, nc9541, nc9542, nc9543, nc9544, nc9545, 
        nc9546, nc9547, nc9548, nc9549, nc9550, nc9551, nc9552, nc9553, 
        nc9554, \A_DOUT_TEMPR103[24] , \A_DOUT_TEMPR103[23] , 
        \A_DOUT_TEMPR103[22] , \A_DOUT_TEMPR103[21] , 
        \A_DOUT_TEMPR103[20] }), .B_DOUT({nc9555, nc9556, nc9557, 
        nc9558, nc9559, nc9560, nc9561, nc9562, nc9563, nc9564, nc9565, 
        nc9566, nc9567, nc9568, nc9569, \B_DOUT_TEMPR103[24] , 
        \B_DOUT_TEMPR103[23] , \B_DOUT_TEMPR103[22] , 
        \B_DOUT_TEMPR103[21] , \B_DOUT_TEMPR103[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[103][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1122 (.A(\B_DOUT_TEMPR16[4] ), .B(\B_DOUT_TEMPR17[4] ), .C(
        \B_DOUT_TEMPR18[4] ), .D(\B_DOUT_TEMPR19[4] ), .Y(OR4_1122_Y));
    OR4 OR4_204 (.A(\B_DOUT_TEMPR52[0] ), .B(\B_DOUT_TEMPR53[0] ), .C(
        \B_DOUT_TEMPR54[0] ), .D(\B_DOUT_TEMPR55[0] ), .Y(OR4_204_Y));
    OR4 OR4_2599 (.A(OR4_345_Y), .B(OR4_2885_Y), .C(OR4_1320_Y), .D(
        OR4_2889_Y), .Y(OR4_2599_Y));
    OR4 OR4_2356 (.A(\B_DOUT_TEMPR60[12] ), .B(\B_DOUT_TEMPR61[12] ), 
        .C(\B_DOUT_TEMPR62[12] ), .D(\B_DOUT_TEMPR63[12] ), .Y(
        OR4_2356_Y));
    OR4 OR4_856 (.A(\B_DOUT_TEMPR111[13] ), .B(\B_DOUT_TEMPR112[13] ), 
        .C(\B_DOUT_TEMPR113[13] ), .D(\B_DOUT_TEMPR114[13] ), .Y(
        OR4_856_Y));
    OR4 OR4_1293 (.A(\A_DOUT_TEMPR24[5] ), .B(\A_DOUT_TEMPR25[5] ), .C(
        \A_DOUT_TEMPR26[5] ), .D(\A_DOUT_TEMPR27[5] ), .Y(OR4_1293_Y));
    OR4 OR4_2778 (.A(\B_DOUT_TEMPR107[26] ), .B(\B_DOUT_TEMPR108[26] ), 
        .C(\B_DOUT_TEMPR109[26] ), .D(\B_DOUT_TEMPR110[26] ), .Y(
        OR4_2778_Y));
    OR4 OR4_1702 (.A(\B_DOUT_TEMPR16[33] ), .B(\B_DOUT_TEMPR17[33] ), 
        .C(\B_DOUT_TEMPR18[33] ), .D(\B_DOUT_TEMPR19[33] ), .Y(
        OR4_1702_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%21%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R21C3 (
        .A_DOUT({nc9570, nc9571, nc9572, nc9573, nc9574, nc9575, 
        nc9576, nc9577, nc9578, nc9579, nc9580, nc9581, nc9582, nc9583, 
        nc9584, \A_DOUT_TEMPR21[19] , \A_DOUT_TEMPR21[18] , 
        \A_DOUT_TEMPR21[17] , \A_DOUT_TEMPR21[16] , 
        \A_DOUT_TEMPR21[15] }), .B_DOUT({nc9585, nc9586, nc9587, 
        nc9588, nc9589, nc9590, nc9591, nc9592, nc9593, nc9594, nc9595, 
        nc9596, nc9597, nc9598, nc9599, \B_DOUT_TEMPR21[19] , 
        \B_DOUT_TEMPR21[18] , \B_DOUT_TEMPR21[17] , 
        \B_DOUT_TEMPR21[16] , \B_DOUT_TEMPR21[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[21][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1964 (.A(\A_DOUT_TEMPR32[16] ), .B(\A_DOUT_TEMPR33[16] ), 
        .C(\A_DOUT_TEMPR34[16] ), .D(\A_DOUT_TEMPR35[16] ), .Y(
        OR4_1964_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%83%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R83C5 (
        .A_DOUT({nc9600, nc9601, nc9602, nc9603, nc9604, nc9605, 
        nc9606, nc9607, nc9608, nc9609, nc9610, nc9611, nc9612, nc9613, 
        nc9614, \A_DOUT_TEMPR83[29] , \A_DOUT_TEMPR83[28] , 
        \A_DOUT_TEMPR83[27] , \A_DOUT_TEMPR83[26] , 
        \A_DOUT_TEMPR83[25] }), .B_DOUT({nc9615, nc9616, nc9617, 
        nc9618, nc9619, nc9620, nc9621, nc9622, nc9623, nc9624, nc9625, 
        nc9626, nc9627, nc9628, nc9629, \B_DOUT_TEMPR83[29] , 
        \B_DOUT_TEMPR83[28] , \B_DOUT_TEMPR83[27] , 
        \B_DOUT_TEMPR83[26] , \B_DOUT_TEMPR83[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[83][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_700 (.A(\A_DOUT_TEMPR64[28] ), .B(\A_DOUT_TEMPR65[28] ), 
        .C(\A_DOUT_TEMPR66[28] ), .D(\A_DOUT_TEMPR67[28] ), .Y(
        OR4_700_Y));
    OR4 OR4_350 (.A(OR4_2987_Y), .B(OR4_1998_Y), .C(OR4_2180_Y), .D(
        OR4_2011_Y), .Y(OR4_350_Y));
    OR4 OR4_18 (.A(OR4_183_Y), .B(OR4_1128_Y), .C(OR4_749_Y), .D(
        OR4_2234_Y), .Y(OR4_18_Y));
    OR4 OR4_789 (.A(\A_DOUT_TEMPR4[3] ), .B(\A_DOUT_TEMPR5[3] ), .C(
        \A_DOUT_TEMPR6[3] ), .D(\A_DOUT_TEMPR7[3] ), .Y(OR4_789_Y));
    OR4 OR4_2392 (.A(\B_DOUT_TEMPR44[34] ), .B(\B_DOUT_TEMPR45[34] ), 
        .C(\B_DOUT_TEMPR46[34] ), .D(\B_DOUT_TEMPR47[34] ), .Y(
        OR4_2392_Y));
    OR4 OR4_1966 (.A(\B_DOUT_TEMPR36[30] ), .B(\B_DOUT_TEMPR37[30] ), 
        .C(\B_DOUT_TEMPR38[30] ), .D(\B_DOUT_TEMPR39[30] ), .Y(
        OR4_1966_Y));
    OR4 OR4_2104 (.A(\A_DOUT_TEMPR20[30] ), .B(\A_DOUT_TEMPR21[30] ), 
        .C(\A_DOUT_TEMPR22[30] ), .D(\A_DOUT_TEMPR23[30] ), .Y(
        OR4_2104_Y));
    OR4 OR4_685 (.A(\A_DOUT_TEMPR0[37] ), .B(\A_DOUT_TEMPR1[37] ), .C(
        \A_DOUT_TEMPR2[37] ), .D(\A_DOUT_TEMPR3[37] ), .Y(OR4_685_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%2%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R2C5 (
        .A_DOUT({nc9630, nc9631, nc9632, nc9633, nc9634, nc9635, 
        nc9636, nc9637, nc9638, nc9639, nc9640, nc9641, nc9642, nc9643, 
        nc9644, \A_DOUT_TEMPR2[29] , \A_DOUT_TEMPR2[28] , 
        \A_DOUT_TEMPR2[27] , \A_DOUT_TEMPR2[26] , \A_DOUT_TEMPR2[25] })
        , .B_DOUT({nc9645, nc9646, nc9647, nc9648, nc9649, nc9650, 
        nc9651, nc9652, nc9653, nc9654, nc9655, nc9656, nc9657, nc9658, 
        nc9659, \B_DOUT_TEMPR2[29] , \B_DOUT_TEMPR2[28] , 
        \B_DOUT_TEMPR2[27] , \B_DOUT_TEMPR2[26] , \B_DOUT_TEMPR2[25] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[2][5] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], \BLKX0[0] }), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[29], A_DIN[28], A_DIN[27], 
        A_DIN[26], A_DIN[25]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2089 (.A(\A_DOUT_TEMPR75[6] ), .B(\A_DOUT_TEMPR76[6] ), .C(
        \A_DOUT_TEMPR77[6] ), .D(\A_DOUT_TEMPR78[6] ), .Y(OR4_2089_Y));
    OR4 OR4_1583 (.A(\B_DOUT_TEMPR87[8] ), .B(\B_DOUT_TEMPR88[8] ), .C(
        \B_DOUT_TEMPR89[8] ), .D(\B_DOUT_TEMPR90[8] ), .Y(OR4_1583_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%41%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R41C5 (
        .A_DOUT({nc9660, nc9661, nc9662, nc9663, nc9664, nc9665, 
        nc9666, nc9667, nc9668, nc9669, nc9670, nc9671, nc9672, nc9673, 
        nc9674, \A_DOUT_TEMPR41[29] , \A_DOUT_TEMPR41[28] , 
        \A_DOUT_TEMPR41[27] , \A_DOUT_TEMPR41[26] , 
        \A_DOUT_TEMPR41[25] }), .B_DOUT({nc9675, nc9676, nc9677, 
        nc9678, nc9679, nc9680, nc9681, nc9682, nc9683, nc9684, nc9685, 
        nc9686, nc9687, nc9688, nc9689, \B_DOUT_TEMPR41[29] , 
        \B_DOUT_TEMPR41[28] , \B_DOUT_TEMPR41[27] , 
        \B_DOUT_TEMPR41[26] , \B_DOUT_TEMPR41[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[41][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[7]  (.A(OR4_2835_Y), .B(OR4_2868_Y), .C(OR4_55_Y), 
        .D(OR4_1626_Y), .Y(B_DOUT[7]));
    OR4 OR4_1412 (.A(OR4_365_Y), .B(OR4_672_Y), .C(OR4_292_Y), .D(
        OR4_692_Y), .Y(OR4_1412_Y));
    OR4 OR4_1758 (.A(OR4_2099_Y), .B(OR4_630_Y), .C(OR4_1453_Y), .D(
        OR4_488_Y), .Y(OR4_1758_Y));
    OR4 OR4_262 (.A(\A_DOUT_TEMPR52[14] ), .B(\A_DOUT_TEMPR53[14] ), 
        .C(\A_DOUT_TEMPR54[14] ), .D(\A_DOUT_TEMPR55[14] ), .Y(
        OR4_262_Y));
    OR4 OR4_194 (.A(OR4_2082_Y), .B(OR4_2204_Y), .C(OR4_1414_Y), .D(
        OR4_334_Y), .Y(OR4_194_Y));
    OR4 OR4_394 (.A(OR4_866_Y), .B(OR4_2912_Y), .C(OR4_542_Y), .D(
        OR4_848_Y), .Y(OR4_394_Y));
    OR4 OR4_289 (.A(\A_DOUT_TEMPR83[6] ), .B(\A_DOUT_TEMPR84[6] ), .C(
        \A_DOUT_TEMPR85[6] ), .D(\A_DOUT_TEMPR86[6] ), .Y(OR4_289_Y));
    OR4 OR4_1240 (.A(\B_DOUT_TEMPR8[38] ), .B(\B_DOUT_TEMPR9[38] ), .C(
        \B_DOUT_TEMPR10[38] ), .D(\B_DOUT_TEMPR11[38] ), .Y(OR4_1240_Y)
        );
    OR4 OR4_2589 (.A(\A_DOUT_TEMPR99[15] ), .B(\A_DOUT_TEMPR100[15] ), 
        .C(\A_DOUT_TEMPR101[15] ), .D(\A_DOUT_TEMPR102[15] ), .Y(
        OR4_2589_Y));
    OR4 OR4_1418 (.A(\A_DOUT_TEMPR115[28] ), .B(\A_DOUT_TEMPR116[28] ), 
        .C(\A_DOUT_TEMPR117[28] ), .D(\A_DOUT_TEMPR118[28] ), .Y(
        OR4_1418_Y));
    OR4 OR4_1183 (.A(\B_DOUT_TEMPR8[1] ), .B(\B_DOUT_TEMPR9[1] ), .C(
        \B_DOUT_TEMPR10[1] ), .D(\B_DOUT_TEMPR11[1] ), .Y(OR4_1183_Y));
    OR4 OR4_1602 (.A(\B_DOUT_TEMPR0[26] ), .B(\B_DOUT_TEMPR1[26] ), .C(
        \B_DOUT_TEMPR2[26] ), .D(\B_DOUT_TEMPR3[26] ), .Y(OR4_1602_Y));
    OR4 OR4_2138 (.A(\B_DOUT_TEMPR44[37] ), .B(\B_DOUT_TEMPR45[37] ), 
        .C(\B_DOUT_TEMPR46[37] ), .D(\B_DOUT_TEMPR47[37] ), .Y(
        OR4_2138_Y));
    OR4 OR4_783 (.A(OR4_1378_Y), .B(OR4_2706_Y), .C(OR4_2317_Y), .D(
        OR4_337_Y), .Y(OR4_783_Y));
    OR4 OR4_1082 (.A(\A_DOUT_TEMPR40[7] ), .B(\A_DOUT_TEMPR41[7] ), .C(
        \A_DOUT_TEMPR42[7] ), .D(\A_DOUT_TEMPR43[7] ), .Y(OR4_1082_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%20%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R20C2 (
        .A_DOUT({nc9690, nc9691, nc9692, nc9693, nc9694, nc9695, 
        nc9696, nc9697, nc9698, nc9699, nc9700, nc9701, nc9702, nc9703, 
        nc9704, \A_DOUT_TEMPR20[14] , \A_DOUT_TEMPR20[13] , 
        \A_DOUT_TEMPR20[12] , \A_DOUT_TEMPR20[11] , 
        \A_DOUT_TEMPR20[10] }), .B_DOUT({nc9705, nc9706, nc9707, 
        nc9708, nc9709, nc9710, nc9711, nc9712, nc9713, nc9714, nc9715, 
        nc9716, nc9717, nc9718, nc9719, \B_DOUT_TEMPR20[14] , 
        \B_DOUT_TEMPR20[13] , \B_DOUT_TEMPR20[12] , 
        \B_DOUT_TEMPR20[11] , \B_DOUT_TEMPR20[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[20][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1138 (.A(\B_DOUT_TEMPR111[27] ), .B(\B_DOUT_TEMPR112[27] ), 
        .C(\B_DOUT_TEMPR113[27] ), .D(\B_DOUT_TEMPR114[27] ), .Y(
        OR4_1138_Y));
    OR4 OR4_1902 (.A(\B_DOUT_TEMPR12[22] ), .B(\B_DOUT_TEMPR13[22] ), 
        .C(\B_DOUT_TEMPR14[22] ), .D(\B_DOUT_TEMPR15[22] ), .Y(
        OR4_1902_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%86%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R86C4 (
        .A_DOUT({nc9720, nc9721, nc9722, nc9723, nc9724, nc9725, 
        nc9726, nc9727, nc9728, nc9729, nc9730, nc9731, nc9732, nc9733, 
        nc9734, \A_DOUT_TEMPR86[24] , \A_DOUT_TEMPR86[23] , 
        \A_DOUT_TEMPR86[22] , \A_DOUT_TEMPR86[21] , 
        \A_DOUT_TEMPR86[20] }), .B_DOUT({nc9735, nc9736, nc9737, 
        nc9738, nc9739, nc9740, nc9741, nc9742, nc9743, nc9744, nc9745, 
        nc9746, nc9747, nc9748, nc9749, \B_DOUT_TEMPR86[24] , 
        \B_DOUT_TEMPR86[23] , \B_DOUT_TEMPR86[22] , 
        \B_DOUT_TEMPR86[21] , \B_DOUT_TEMPR86[20] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[86][4] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[24], A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[24], 
        B_DIN[23], B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_240 (.A(OR4_1521_Y), .B(OR4_2739_Y), .C(OR2_23_Y), .D(
        \A_DOUT_TEMPR74[16] ), .Y(OR4_240_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%3%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R3C5 (
        .A_DOUT({nc9750, nc9751, nc9752, nc9753, nc9754, nc9755, 
        nc9756, nc9757, nc9758, nc9759, nc9760, nc9761, nc9762, nc9763, 
        nc9764, \A_DOUT_TEMPR3[29] , \A_DOUT_TEMPR3[28] , 
        \A_DOUT_TEMPR3[27] , \A_DOUT_TEMPR3[26] , \A_DOUT_TEMPR3[25] })
        , .B_DOUT({nc9765, nc9766, nc9767, nc9768, nc9769, nc9770, 
        nc9771, nc9772, nc9773, nc9774, nc9775, nc9776, nc9777, nc9778, 
        nc9779, \B_DOUT_TEMPR3[29] , \B_DOUT_TEMPR3[28] , 
        \B_DOUT_TEMPR3[27] , \B_DOUT_TEMPR3[26] , \B_DOUT_TEMPR3[25] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[3][5] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], A_ADDR[12]}), .A_CLK(
        A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, A_DIN[29], A_DIN[28], A_DIN[27], 
        A_DIN[26], A_DIN[25]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2382 (.A(\A_DOUT_TEMPR0[19] ), .B(\A_DOUT_TEMPR1[19] ), .C(
        \A_DOUT_TEMPR2[19] ), .D(\A_DOUT_TEMPR3[19] ), .Y(OR4_2382_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%54%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R54C0 (
        .A_DOUT({nc9780, nc9781, nc9782, nc9783, nc9784, nc9785, 
        nc9786, nc9787, nc9788, nc9789, nc9790, nc9791, nc9792, nc9793, 
        nc9794, \A_DOUT_TEMPR54[4] , \A_DOUT_TEMPR54[3] , 
        \A_DOUT_TEMPR54[2] , \A_DOUT_TEMPR54[1] , \A_DOUT_TEMPR54[0] })
        , .B_DOUT({nc9795, nc9796, nc9797, nc9798, nc9799, nc9800, 
        nc9801, nc9802, nc9803, nc9804, nc9805, nc9806, nc9807, nc9808, 
        nc9809, \B_DOUT_TEMPR54[4] , \B_DOUT_TEMPR54[3] , 
        \B_DOUT_TEMPR54[2] , \B_DOUT_TEMPR54[1] , \B_DOUT_TEMPR54[0] })
        , .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(
        \ACCESS_BUSY[54][0] ), .A_ADDR({A_ADDR[11], A_ADDR[10], 
        A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], A_ADDR[5], 
        A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, 
        GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], \BLKX0[0] }), 
        .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, A_DIN[4], A_DIN[3], 
        A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, 
        \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), 
        .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%17%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R17C5 (
        .A_DOUT({nc9810, nc9811, nc9812, nc9813, nc9814, nc9815, 
        nc9816, nc9817, nc9818, nc9819, nc9820, nc9821, nc9822, nc9823, 
        nc9824, \A_DOUT_TEMPR17[29] , \A_DOUT_TEMPR17[28] , 
        \A_DOUT_TEMPR17[27] , \A_DOUT_TEMPR17[26] , 
        \A_DOUT_TEMPR17[25] }), .B_DOUT({nc9825, nc9826, nc9827, 
        nc9828, nc9829, nc9830, nc9831, nc9832, nc9833, nc9834, nc9835, 
        nc9836, nc9837, nc9838, nc9839, \B_DOUT_TEMPR17[29] , 
        \B_DOUT_TEMPR17[28] , \B_DOUT_TEMPR17[27] , 
        \B_DOUT_TEMPR17[26] , \B_DOUT_TEMPR17[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[17][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[0]  (.A(OR4_1635_Y), .B(OR4_29_Y), .C(OR4_1087_Y), 
        .D(OR4_902_Y), .Y(A_DOUT[0]));
    OR4 OR4_640 (.A(\A_DOUT_TEMPR68[15] ), .B(\A_DOUT_TEMPR69[15] ), 
        .C(\A_DOUT_TEMPR70[15] ), .D(\A_DOUT_TEMPR71[15] ), .Y(
        OR4_640_Y));
    OR4 OR4_2833 (.A(\A_DOUT_TEMPR24[9] ), .B(\A_DOUT_TEMPR25[9] ), .C(
        \A_DOUT_TEMPR26[9] ), .D(\A_DOUT_TEMPR27[9] ), .Y(OR4_2833_Y));
    OR4 OR4_2805 (.A(\A_DOUT_TEMPR99[26] ), .B(\A_DOUT_TEMPR100[26] ), 
        .C(\A_DOUT_TEMPR101[26] ), .D(\A_DOUT_TEMPR102[26] ), .Y(
        OR4_2805_Y));
    OR4 OR4_2595 (.A(\A_DOUT_TEMPR4[15] ), .B(\A_DOUT_TEMPR5[15] ), .C(
        \A_DOUT_TEMPR6[15] ), .D(\A_DOUT_TEMPR7[15] ), .Y(OR4_2595_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%99%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R99C3 (
        .A_DOUT({nc9840, nc9841, nc9842, nc9843, nc9844, nc9845, 
        nc9846, nc9847, nc9848, nc9849, nc9850, nc9851, nc9852, nc9853, 
        nc9854, \A_DOUT_TEMPR99[19] , \A_DOUT_TEMPR99[18] , 
        \A_DOUT_TEMPR99[17] , \A_DOUT_TEMPR99[16] , 
        \A_DOUT_TEMPR99[15] }), .B_DOUT({nc9855, nc9856, nc9857, 
        nc9858, nc9859, nc9860, nc9861, nc9862, nc9863, nc9864, nc9865, 
        nc9866, nc9867, nc9868, nc9869, \B_DOUT_TEMPR99[19] , 
        \B_DOUT_TEMPR99[18] , \B_DOUT_TEMPR99[17] , 
        \B_DOUT_TEMPR99[16] , \B_DOUT_TEMPR99[15] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[99][3] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[19], A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[19], 
        B_DIN[18], B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1510 (.A(OR4_1680_Y), .B(OR4_1496_Y), .C(OR4_1443_Y), .D(
        OR4_1544_Y), .Y(OR4_1510_Y));
    OR4 OR4_288 (.A(\A_DOUT_TEMPR8[8] ), .B(\A_DOUT_TEMPR9[8] ), .C(
        \A_DOUT_TEMPR10[8] ), .D(\A_DOUT_TEMPR11[8] ), .Y(OR4_288_Y));
    OR4 OR4_1346 (.A(\B_DOUT_TEMPR103[3] ), .B(\B_DOUT_TEMPR104[3] ), 
        .C(\B_DOUT_TEMPR105[3] ), .D(\B_DOUT_TEMPR106[3] ), .Y(
        OR4_1346_Y));
    OR4 OR4_2452 (.A(\A_DOUT_TEMPR83[7] ), .B(\A_DOUT_TEMPR84[7] ), .C(
        \A_DOUT_TEMPR85[7] ), .D(\A_DOUT_TEMPR86[7] ), .Y(OR4_2452_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%85%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R85C5 (
        .A_DOUT({nc9870, nc9871, nc9872, nc9873, nc9874, nc9875, 
        nc9876, nc9877, nc9878, nc9879, nc9880, nc9881, nc9882, nc9883, 
        nc9884, \A_DOUT_TEMPR85[29] , \A_DOUT_TEMPR85[28] , 
        \A_DOUT_TEMPR85[27] , \A_DOUT_TEMPR85[26] , 
        \A_DOUT_TEMPR85[25] }), .B_DOUT({nc9885, nc9886, nc9887, 
        nc9888, nc9889, nc9890, nc9891, nc9892, nc9893, nc9894, nc9895, 
        nc9896, nc9897, nc9898, nc9899, \B_DOUT_TEMPR85[29] , 
        \B_DOUT_TEMPR85[28] , \B_DOUT_TEMPR85[27] , 
        \B_DOUT_TEMPR85[26] , \B_DOUT_TEMPR85[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[85][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR2 OR2_8 (.A(\A_DOUT_TEMPR72[8] ), .B(\A_DOUT_TEMPR73[8] ), .Y(
        OR2_8_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%67%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R67C2 (
        .A_DOUT({nc9900, nc9901, nc9902, nc9903, nc9904, nc9905, 
        nc9906, nc9907, nc9908, nc9909, nc9910, nc9911, nc9912, nc9913, 
        nc9914, \A_DOUT_TEMPR67[14] , \A_DOUT_TEMPR67[13] , 
        \A_DOUT_TEMPR67[12] , \A_DOUT_TEMPR67[11] , 
        \A_DOUT_TEMPR67[10] }), .B_DOUT({nc9915, nc9916, nc9917, 
        nc9918, nc9919, nc9920, nc9921, nc9922, nc9923, nc9924, nc9925, 
        nc9926, nc9927, nc9928, nc9929, \B_DOUT_TEMPR67[14] , 
        \B_DOUT_TEMPR67[13] , \B_DOUT_TEMPR67[12] , 
        \B_DOUT_TEMPR67[11] , \B_DOUT_TEMPR67[10] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[67][2] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , 
        A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[14], A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], 
        B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[14], 
        B_DIN[13], B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1833 (.A(\A_DOUT_TEMPR28[11] ), .B(\A_DOUT_TEMPR29[11] ), 
        .C(\A_DOUT_TEMPR30[11] ), .D(\A_DOUT_TEMPR31[11] ), .Y(
        OR4_1833_Y));
    OR2 OR2_23 (.A(\A_DOUT_TEMPR72[16] ), .B(\A_DOUT_TEMPR73[16] ), .Y(
        OR2_23_Y));
    OR4 OR4_1079 (.A(OR4_2614_Y), .B(OR4_380_Y), .C(OR2_63_Y), .D(
        \B_DOUT_TEMPR74[29] ), .Y(OR4_1079_Y));
    OR4 OR4_2458 (.A(\A_DOUT_TEMPR32[35] ), .B(\A_DOUT_TEMPR33[35] ), 
        .C(\A_DOUT_TEMPR34[35] ), .D(\A_DOUT_TEMPR35[35] ), .Y(
        OR4_2458_Y));
    OR4 OR4_2739 (.A(\A_DOUT_TEMPR68[16] ), .B(\A_DOUT_TEMPR69[16] ), 
        .C(\A_DOUT_TEMPR70[16] ), .D(\A_DOUT_TEMPR71[16] ), .Y(
        OR4_2739_Y));
    OR4 OR4_2523 (.A(OR4_1522_Y), .B(OR4_2432_Y), .C(OR4_2086_Y), .D(
        OR4_548_Y), .Y(OR4_2523_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%84%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R84C5 (
        .A_DOUT({nc9930, nc9931, nc9932, nc9933, nc9934, nc9935, 
        nc9936, nc9937, nc9938, nc9939, nc9940, nc9941, nc9942, nc9943, 
        nc9944, \A_DOUT_TEMPR84[29] , \A_DOUT_TEMPR84[28] , 
        \A_DOUT_TEMPR84[27] , \A_DOUT_TEMPR84[26] , 
        \A_DOUT_TEMPR84[25] }), .B_DOUT({nc9945, nc9946, nc9947, 
        nc9948, nc9949, nc9950, nc9951, nc9952, nc9953, nc9954, nc9955, 
        nc9956, nc9957, nc9958, nc9959, \B_DOUT_TEMPR84[29] , 
        \B_DOUT_TEMPR84[28] , \B_DOUT_TEMPR84[27] , 
        \B_DOUT_TEMPR84[26] , \B_DOUT_TEMPR84[25] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[84][5] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[29], A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[29], 
        B_DIN[28], B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_2410 (.A(\A_DOUT_TEMPR12[10] ), .B(\A_DOUT_TEMPR13[10] ), 
        .C(\A_DOUT_TEMPR14[10] ), .D(\A_DOUT_TEMPR15[10] ), .Y(
        OR4_2410_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%56%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R56C7 (
        .A_DOUT({nc9960, nc9961, nc9962, nc9963, nc9964, nc9965, 
        nc9966, nc9967, nc9968, nc9969, nc9970, nc9971, nc9972, nc9973, 
        nc9974, \A_DOUT_TEMPR56[39] , \A_DOUT_TEMPR56[38] , 
        \A_DOUT_TEMPR56[37] , \A_DOUT_TEMPR56[36] , 
        \A_DOUT_TEMPR56[35] }), .B_DOUT({nc9975, nc9976, nc9977, 
        nc9978, nc9979, nc9980, nc9981, nc9982, nc9983, nc9984, nc9985, 
        nc9986, nc9987, nc9988, nc9989, \B_DOUT_TEMPR56[39] , 
        \B_DOUT_TEMPR56[38] , \B_DOUT_TEMPR56[37] , 
        \B_DOUT_TEMPR56[36] , \B_DOUT_TEMPR56[35] }), .DB_DETECT(), 
        .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[56][7] ), .A_ADDR({
        A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], 
        A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], 
        A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , 
        \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        A_DIN[39], A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), 
        .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), 
        .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], 
        B_ADDR[10], B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], 
        B_ADDR[5], B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], 
        B_ADDR[0], GND, GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , 
        \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, B_DIN[39], 
        B_DIN[38], B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), 
        .B_WEN({GND, \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(
        VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), 
        .A_WIDTH({GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC)
        , .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(
        VCC), .ECC_BYPASS(GND));
    OR4 OR4_1579 (.A(\B_DOUT_TEMPR52[6] ), .B(\B_DOUT_TEMPR53[6] ), .C(
        \B_DOUT_TEMPR54[6] ), .D(\B_DOUT_TEMPR55[6] ), .Y(OR4_1579_Y));
    OR4 OR4_1739 (.A(\A_DOUT_TEMPR103[34] ), .B(\A_DOUT_TEMPR104[34] ), 
        .C(\A_DOUT_TEMPR105[34] ), .D(\A_DOUT_TEMPR106[34] ), .Y(
        OR4_1739_Y));
    OR4 OR4_2123 (.A(\B_DOUT_TEMPR40[39] ), .B(\B_DOUT_TEMPR41[39] ), 
        .C(\B_DOUT_TEMPR42[39] ), .D(\B_DOUT_TEMPR43[39] ), .Y(
        OR4_2123_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%101%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R101C6 (
        .A_DOUT({nc9990, nc9991, nc9992, nc9993, nc9994, nc9995, 
        nc9996, nc9997, nc9998, nc9999, nc10000, nc10001, nc10002, 
        nc10003, nc10004, \A_DOUT_TEMPR101[34] , \A_DOUT_TEMPR101[33] , 
        \A_DOUT_TEMPR101[32] , \A_DOUT_TEMPR101[31] , 
        \A_DOUT_TEMPR101[30] }), .B_DOUT({nc10005, nc10006, nc10007, 
        nc10008, nc10009, nc10010, nc10011, nc10012, nc10013, nc10014, 
        nc10015, nc10016, nc10017, nc10018, nc10019, 
        \B_DOUT_TEMPR101[34] , \B_DOUT_TEMPR101[33] , 
        \B_DOUT_TEMPR101[32] , \B_DOUT_TEMPR101[31] , 
        \B_DOUT_TEMPR101[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[101][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%57%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R57C6 (
        .A_DOUT({nc10020, nc10021, nc10022, nc10023, nc10024, nc10025, 
        nc10026, nc10027, nc10028, nc10029, nc10030, nc10031, nc10032, 
        nc10033, nc10034, \A_DOUT_TEMPR57[34] , \A_DOUT_TEMPR57[33] , 
        \A_DOUT_TEMPR57[32] , \A_DOUT_TEMPR57[31] , 
        \A_DOUT_TEMPR57[30] }), .B_DOUT({nc10035, nc10036, nc10037, 
        nc10038, nc10039, nc10040, nc10041, nc10042, nc10043, nc10044, 
        nc10045, nc10046, nc10047, nc10048, nc10049, 
        \B_DOUT_TEMPR57[34] , \B_DOUT_TEMPR57[33] , 
        \B_DOUT_TEMPR57[32] , \B_DOUT_TEMPR57[31] , 
        \B_DOUT_TEMPR57[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[57][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2136 (.A(\B_DOUT_TEMPR12[1] ), .B(\B_DOUT_TEMPR13[1] ), .C(
        \B_DOUT_TEMPR14[1] ), .D(\B_DOUT_TEMPR15[1] ), .Y(OR4_2136_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%101%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R101C7 (
        .A_DOUT({nc10050, nc10051, nc10052, nc10053, nc10054, nc10055, 
        nc10056, nc10057, nc10058, nc10059, nc10060, nc10061, nc10062, 
        nc10063, nc10064, \A_DOUT_TEMPR101[39] , \A_DOUT_TEMPR101[38] , 
        \A_DOUT_TEMPR101[37] , \A_DOUT_TEMPR101[36] , 
        \A_DOUT_TEMPR101[35] }), .B_DOUT({nc10065, nc10066, nc10067, 
        nc10068, nc10069, nc10070, nc10071, nc10072, nc10073, nc10074, 
        nc10075, nc10076, nc10077, nc10078, nc10079, 
        \B_DOUT_TEMPR101[39] , \B_DOUT_TEMPR101[38] , 
        \B_DOUT_TEMPR101[37] , \B_DOUT_TEMPR101[36] , 
        \B_DOUT_TEMPR101[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[101][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%97%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R97C3 (
        .A_DOUT({nc10080, nc10081, nc10082, nc10083, nc10084, nc10085, 
        nc10086, nc10087, nc10088, nc10089, nc10090, nc10091, nc10092, 
        nc10093, nc10094, \A_DOUT_TEMPR97[19] , \A_DOUT_TEMPR97[18] , 
        \A_DOUT_TEMPR97[17] , \A_DOUT_TEMPR97[16] , 
        \A_DOUT_TEMPR97[15] }), .B_DOUT({nc10095, nc10096, nc10097, 
        nc10098, nc10099, nc10100, nc10101, nc10102, nc10103, nc10104, 
        nc10105, nc10106, nc10107, nc10108, nc10109, 
        \B_DOUT_TEMPR97[19] , \B_DOUT_TEMPR97[18] , 
        \B_DOUT_TEMPR97[17] , \B_DOUT_TEMPR97[16] , 
        \B_DOUT_TEMPR97[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[97][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2585 (.A(OR4_2941_Y), .B(OR4_1550_Y), .C(OR4_1020_Y), .D(
        OR4_2302_Y), .Y(OR4_2585_Y));
    OR4 OR4_2022 (.A(\B_DOUT_TEMPR79[27] ), .B(\B_DOUT_TEMPR80[27] ), 
        .C(\B_DOUT_TEMPR81[27] ), .D(\B_DOUT_TEMPR82[27] ), .Y(
        OR4_2022_Y));
    OR4 OR4_2538 (.A(\A_DOUT_TEMPR68[21] ), .B(\A_DOUT_TEMPR69[21] ), 
        .C(\A_DOUT_TEMPR70[21] ), .D(\A_DOUT_TEMPR71[21] ), .Y(
        OR4_2538_Y));
    OR4 OR4_254 (.A(\B_DOUT_TEMPR91[25] ), .B(\B_DOUT_TEMPR92[25] ), 
        .C(\B_DOUT_TEMPR93[25] ), .D(\B_DOUT_TEMPR94[25] ), .Y(
        OR4_254_Y));
    OR4 OR4_233 (.A(\B_DOUT_TEMPR20[38] ), .B(\B_DOUT_TEMPR21[38] ), 
        .C(\B_DOUT_TEMPR22[38] ), .D(\B_DOUT_TEMPR23[38] ), .Y(
        OR4_233_Y));
    OR4 OR4_2215 (.A(\A_DOUT_TEMPR83[37] ), .B(\A_DOUT_TEMPR84[37] ), 
        .C(\A_DOUT_TEMPR85[37] ), .D(\A_DOUT_TEMPR86[37] ), .Y(
        OR4_2215_Y));
    OR4 OR4_2550 (.A(OR4_130_Y), .B(OR4_980_Y), .C(OR2_0_Y), .D(
        \A_DOUT_TEMPR74[27] ), .Y(OR4_2550_Y));
    OR4 OR4_1372 (.A(OR4_2246_Y), .B(OR4_2079_Y), .C(OR4_2032_Y), .D(
        OR4_1069_Y), .Y(OR4_1372_Y));
    OR4 OR4_1136 (.A(\B_DOUT_TEMPR107[7] ), .B(\B_DOUT_TEMPR108[7] ), 
        .C(\B_DOUT_TEMPR109[7] ), .D(\B_DOUT_TEMPR110[7] ), .Y(
        OR4_1136_Y));
    OR4 OR4_331 (.A(\B_DOUT_TEMPR99[19] ), .B(\B_DOUT_TEMPR100[19] ), 
        .C(\B_DOUT_TEMPR101[19] ), .D(\B_DOUT_TEMPR102[19] ), .Y(
        OR4_331_Y));
    OR4 OR4_1229 (.A(\B_DOUT_TEMPR24[2] ), .B(\B_DOUT_TEMPR25[2] ), .C(
        \B_DOUT_TEMPR26[2] ), .D(\B_DOUT_TEMPR27[2] ), .Y(OR4_1229_Y));
    OR4 OR4_835 (.A(\A_DOUT_TEMPR24[13] ), .B(\A_DOUT_TEMPR25[13] ), 
        .C(\A_DOUT_TEMPR26[13] ), .D(\A_DOUT_TEMPR27[13] ), .Y(
        OR4_835_Y));
    OR4 OR4_1538 (.A(\A_DOUT_TEMPR107[24] ), .B(\A_DOUT_TEMPR108[24] ), 
        .C(\A_DOUT_TEMPR109[24] ), .D(\A_DOUT_TEMPR110[24] ), .Y(
        OR4_1538_Y));
    OR4 OR4_28 (.A(\B_DOUT_TEMPR32[17] ), .B(\B_DOUT_TEMPR33[17] ), .C(
        \B_DOUT_TEMPR34[17] ), .D(\B_DOUT_TEMPR35[17] ), .Y(OR4_28_Y));
    OR4 OR4_133 (.A(\A_DOUT_TEMPR16[28] ), .B(\A_DOUT_TEMPR17[28] ), 
        .C(\A_DOUT_TEMPR18[28] ), .D(\A_DOUT_TEMPR19[28] ), .Y(
        OR4_133_Y));
    OR4 OR4_2998 (.A(\A_DOUT_TEMPR60[28] ), .B(\A_DOUT_TEMPR61[28] ), 
        .C(\A_DOUT_TEMPR62[28] ), .D(\A_DOUT_TEMPR63[28] ), .Y(
        OR4_2998_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%15%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R15C7 (
        .A_DOUT({nc10110, nc10111, nc10112, nc10113, nc10114, nc10115, 
        nc10116, nc10117, nc10118, nc10119, nc10120, nc10121, nc10122, 
        nc10123, nc10124, \A_DOUT_TEMPR15[39] , \A_DOUT_TEMPR15[38] , 
        \A_DOUT_TEMPR15[37] , \A_DOUT_TEMPR15[36] , 
        \A_DOUT_TEMPR15[35] }), .B_DOUT({nc10125, nc10126, nc10127, 
        nc10128, nc10129, nc10130, nc10131, nc10132, nc10133, nc10134, 
        nc10135, nc10136, nc10137, nc10138, nc10139, 
        \B_DOUT_TEMPR15[39] , \B_DOUT_TEMPR15[38] , 
        \B_DOUT_TEMPR15[37] , \B_DOUT_TEMPR15[36] , 
        \B_DOUT_TEMPR15[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%52%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R52C4 (
        .A_DOUT({nc10140, nc10141, nc10142, nc10143, nc10144, nc10145, 
        nc10146, nc10147, nc10148, nc10149, nc10150, nc10151, nc10152, 
        nc10153, nc10154, \A_DOUT_TEMPR52[24] , \A_DOUT_TEMPR52[23] , 
        \A_DOUT_TEMPR52[22] , \A_DOUT_TEMPR52[21] , 
        \A_DOUT_TEMPR52[20] }), .B_DOUT({nc10155, nc10156, nc10157, 
        nc10158, nc10159, nc10160, nc10161, nc10162, nc10163, nc10164, 
        nc10165, nc10166, nc10167, nc10168, nc10169, 
        \B_DOUT_TEMPR52[24] , \B_DOUT_TEMPR52[23] , 
        \B_DOUT_TEMPR52[22] , \B_DOUT_TEMPR52[21] , 
        \B_DOUT_TEMPR52[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[52][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_750 (.A(\A_DOUT_TEMPR99[22] ), .B(\A_DOUT_TEMPR100[22] ), 
        .C(\A_DOUT_TEMPR101[22] ), .D(\A_DOUT_TEMPR102[22] ), .Y(
        OR4_750_Y));
    OR4 OR4_187 (.A(\A_DOUT_TEMPR79[21] ), .B(\A_DOUT_TEMPR80[21] ), 
        .C(\A_DOUT_TEMPR81[21] ), .D(\A_DOUT_TEMPR82[21] ), .Y(
        OR4_187_Y));
    OR4 OR4_896 (.A(OR4_1033_Y), .B(OR4_1996_Y), .C(OR4_2691_Y), .D(
        OR4_1318_Y), .Y(OR4_896_Y));
    OR4 OR4_916 (.A(\B_DOUT_TEMPR75[9] ), .B(\B_DOUT_TEMPR76[9] ), .C(
        \B_DOUT_TEMPR77[9] ), .D(\B_DOUT_TEMPR78[9] ), .Y(OR4_916_Y));
    OR4 OR4_1915 (.A(\A_DOUT_TEMPR79[4] ), .B(\A_DOUT_TEMPR80[4] ), .C(
        \A_DOUT_TEMPR81[4] ), .D(\A_DOUT_TEMPR82[4] ), .Y(OR4_1915_Y));
    OR4 \OR4_B_DOUT[9]  (.A(OR4_1380_Y), .B(OR4_16_Y), .C(OR4_2946_Y), 
        .D(OR4_1458_Y), .Y(B_DOUT[9]));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[28]  (.A(CFG3_4_Y), .B(
        CFG3_18_Y), .Y(\BLKX2[28] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%34%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R34C0 (
        .A_DOUT({nc10170, nc10171, nc10172, nc10173, nc10174, nc10175, 
        nc10176, nc10177, nc10178, nc10179, nc10180, nc10181, nc10182, 
        nc10183, nc10184, \A_DOUT_TEMPR34[4] , \A_DOUT_TEMPR34[3] , 
        \A_DOUT_TEMPR34[2] , \A_DOUT_TEMPR34[1] , \A_DOUT_TEMPR34[0] })
        , .B_DOUT({nc10185, nc10186, nc10187, nc10188, nc10189, 
        nc10190, nc10191, nc10192, nc10193, nc10194, nc10195, nc10196, 
        nc10197, nc10198, nc10199, \B_DOUT_TEMPR34[4] , 
        \B_DOUT_TEMPR34[3] , \B_DOUT_TEMPR34[2] , \B_DOUT_TEMPR34[1] , 
        \B_DOUT_TEMPR34[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[34][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_390 (.A(\B_DOUT_TEMPR107[29] ), .B(\B_DOUT_TEMPR108[29] ), 
        .C(\B_DOUT_TEMPR109[29] ), .D(\B_DOUT_TEMPR110[29] ), .Y(
        OR4_390_Y));
    OR4 OR4_1409 (.A(\B_DOUT_TEMPR99[30] ), .B(\B_DOUT_TEMPR100[30] ), 
        .C(\B_DOUT_TEMPR101[30] ), .D(\B_DOUT_TEMPR102[30] ), .Y(
        OR4_1409_Y));
    OR4 OR4_1619 (.A(\B_DOUT_TEMPR95[6] ), .B(\B_DOUT_TEMPR96[6] ), .C(
        \B_DOUT_TEMPR97[6] ), .D(\B_DOUT_TEMPR98[6] ), .Y(OR4_1619_Y));
    OR4 OR4_1442 (.A(\A_DOUT_TEMPR52[18] ), .B(\A_DOUT_TEMPR53[18] ), 
        .C(\A_DOUT_TEMPR54[18] ), .D(\A_DOUT_TEMPR55[18] ), .Y(
        OR4_1442_Y));
    CFG3 #( .INIT(8'h40) )  CFG3_23 (.A(A_ADDR[16]), .B(A_ADDR[15]), 
        .C(A_ADDR[14]), .Y(CFG3_23_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%8%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R8C6 (
        .A_DOUT({nc10200, nc10201, nc10202, nc10203, nc10204, nc10205, 
        nc10206, nc10207, nc10208, nc10209, nc10210, nc10211, nc10212, 
        nc10213, nc10214, \A_DOUT_TEMPR8[34] , \A_DOUT_TEMPR8[33] , 
        \A_DOUT_TEMPR8[32] , \A_DOUT_TEMPR8[31] , \A_DOUT_TEMPR8[30] })
        , .B_DOUT({nc10215, nc10216, nc10217, nc10218, nc10219, 
        nc10220, nc10221, nc10222, nc10223, nc10224, nc10225, nc10226, 
        nc10227, nc10228, nc10229, \B_DOUT_TEMPR8[34] , 
        \B_DOUT_TEMPR8[33] , \B_DOUT_TEMPR8[32] , \B_DOUT_TEMPR8[31] , 
        \B_DOUT_TEMPR8[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1448 (.A(OR4_797_Y), .B(OR4_1729_Y), .C(OR4_2426_Y), .D(
        OR4_2756_Y), .Y(OR4_1448_Y));
    OR4 OR4_2988 (.A(OR4_1660_Y), .B(OR4_123_Y), .C(OR4_709_Y), .D(
        OR4_525_Y), .Y(OR4_2988_Y));
    OR4 OR4_1575 (.A(OR4_1880_Y), .B(OR4_1365_Y), .C(OR4_2697_Y), .D(
        OR4_573_Y), .Y(OR4_1575_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[12]  (.A(CFG3_4_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[12] ));
    OR4 OR4_732 (.A(\B_DOUT_TEMPR95[22] ), .B(\B_DOUT_TEMPR96[22] ), 
        .C(\B_DOUT_TEMPR97[22] ), .D(\B_DOUT_TEMPR98[22] ), .Y(
        OR4_732_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[11]  (.A(CFG3_23_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[11] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%36%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R36C7 (
        .A_DOUT({nc10230, nc10231, nc10232, nc10233, nc10234, nc10235, 
        nc10236, nc10237, nc10238, nc10239, nc10240, nc10241, nc10242, 
        nc10243, nc10244, \A_DOUT_TEMPR36[39] , \A_DOUT_TEMPR36[38] , 
        \A_DOUT_TEMPR36[37] , \A_DOUT_TEMPR36[36] , 
        \A_DOUT_TEMPR36[35] }), .B_DOUT({nc10245, nc10246, nc10247, 
        nc10248, nc10249, nc10250, nc10251, nc10252, nc10253, nc10254, 
        nc10255, nc10256, nc10257, nc10258, nc10259, 
        \B_DOUT_TEMPR36[39] , \B_DOUT_TEMPR36[38] , 
        \B_DOUT_TEMPR36[37] , \B_DOUT_TEMPR36[36] , 
        \B_DOUT_TEMPR36[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%24%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R24C6 (
        .A_DOUT({nc10260, nc10261, nc10262, nc10263, nc10264, nc10265, 
        nc10266, nc10267, nc10268, nc10269, nc10270, nc10271, nc10272, 
        nc10273, nc10274, \A_DOUT_TEMPR24[34] , \A_DOUT_TEMPR24[33] , 
        \A_DOUT_TEMPR24[32] , \A_DOUT_TEMPR24[31] , 
        \A_DOUT_TEMPR24[30] }), .B_DOUT({nc10275, nc10276, nc10277, 
        nc10278, nc10279, nc10280, nc10281, nc10282, nc10283, nc10284, 
        nc10285, nc10286, nc10287, nc10288, nc10289, 
        \B_DOUT_TEMPR24[34] , \B_DOUT_TEMPR24[33] , 
        \B_DOUT_TEMPR24[32] , \B_DOUT_TEMPR24[31] , 
        \B_DOUT_TEMPR24[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_336 (.A(\B_DOUT_TEMPR115[31] ), .B(\B_DOUT_TEMPR116[31] ), 
        .C(\B_DOUT_TEMPR117[31] ), .D(\B_DOUT_TEMPR118[31] ), .Y(
        OR4_336_Y));
    OR4 OR4_2179 (.A(\B_DOUT_TEMPR24[6] ), .B(\B_DOUT_TEMPR25[6] ), .C(
        \B_DOUT_TEMPR26[6] ), .D(\B_DOUT_TEMPR27[6] ), .Y(OR4_2179_Y));
    OR4 OR4_2955 (.A(\A_DOUT_TEMPR56[22] ), .B(\A_DOUT_TEMPR57[22] ), 
        .C(\A_DOUT_TEMPR58[22] ), .D(\A_DOUT_TEMPR59[22] ), .Y(
        OR4_2955_Y));
    OR4 OR4_2197 (.A(\A_DOUT_TEMPR0[8] ), .B(\A_DOUT_TEMPR1[8] ), .C(
        \A_DOUT_TEMPR2[8] ), .D(\A_DOUT_TEMPR3[8] ), .Y(OR4_2197_Y));
    OR4 OR4_2694 (.A(\A_DOUT_TEMPR20[33] ), .B(\A_DOUT_TEMPR21[33] ), 
        .C(\A_DOUT_TEMPR22[33] ), .D(\A_DOUT_TEMPR23[33] ), .Y(
        OR4_2694_Y));
    OR4 OR4_176 (.A(\B_DOUT_TEMPR44[17] ), .B(\B_DOUT_TEMPR45[17] ), 
        .C(\B_DOUT_TEMPR46[17] ), .D(\B_DOUT_TEMPR47[17] ), .Y(
        OR4_176_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_3 (.A(VCC), .B(A_ADDR[18]), .C(
        A_ADDR[17]), .Y(CFG3_3_Y));
    OR4 OR4_1300 (.A(\A_DOUT_TEMPR107[12] ), .B(\A_DOUT_TEMPR108[12] ), 
        .C(\A_DOUT_TEMPR109[12] ), .D(\A_DOUT_TEMPR110[12] ), .Y(
        OR4_1300_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%102%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R102C5 (
        .A_DOUT({nc10290, nc10291, nc10292, nc10293, nc10294, nc10295, 
        nc10296, nc10297, nc10298, nc10299, nc10300, nc10301, nc10302, 
        nc10303, nc10304, \A_DOUT_TEMPR102[29] , \A_DOUT_TEMPR102[28] , 
        \A_DOUT_TEMPR102[27] , \A_DOUT_TEMPR102[26] , 
        \A_DOUT_TEMPR102[25] }), .B_DOUT({nc10305, nc10306, nc10307, 
        nc10308, nc10309, nc10310, nc10311, nc10312, nc10313, nc10314, 
        nc10315, nc10316, nc10317, nc10318, nc10319, 
        \B_DOUT_TEMPR102[29] , \B_DOUT_TEMPR102[28] , 
        \B_DOUT_TEMPR102[27] , \B_DOUT_TEMPR102[26] , 
        \B_DOUT_TEMPR102[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[102][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%37%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R37C6 (
        .A_DOUT({nc10320, nc10321, nc10322, nc10323, nc10324, nc10325, 
        nc10326, nc10327, nc10328, nc10329, nc10330, nc10331, nc10332, 
        nc10333, nc10334, \A_DOUT_TEMPR37[34] , \A_DOUT_TEMPR37[33] , 
        \A_DOUT_TEMPR37[32] , \A_DOUT_TEMPR37[31] , 
        \A_DOUT_TEMPR37[30] }), .B_DOUT({nc10335, nc10336, nc10337, 
        nc10338, nc10339, nc10340, nc10341, nc10342, nc10343, nc10344, 
        nc10345, nc10346, nc10347, nc10348, nc10349, 
        \B_DOUT_TEMPR37[34] , \B_DOUT_TEMPR37[33] , 
        \B_DOUT_TEMPR37[32] , \B_DOUT_TEMPR37[31] , 
        \B_DOUT_TEMPR37[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[37][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1407 (.A(OR4_576_Y), .B(OR4_1514_Y), .C(OR4_317_Y), .D(
        OR4_2419_Y), .Y(OR4_1407_Y));
    OR4 OR4_2069 (.A(OR4_1753_Y), .B(OR4_2688_Y), .C(OR4_2305_Y), .D(
        OR4_773_Y), .Y(OR4_2069_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%88%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R88C4 (
        .A_DOUT({nc10350, nc10351, nc10352, nc10353, nc10354, nc10355, 
        nc10356, nc10357, nc10358, nc10359, nc10360, nc10361, nc10362, 
        nc10363, nc10364, \A_DOUT_TEMPR88[24] , \A_DOUT_TEMPR88[23] , 
        \A_DOUT_TEMPR88[22] , \A_DOUT_TEMPR88[21] , 
        \A_DOUT_TEMPR88[20] }), .B_DOUT({nc10365, nc10366, nc10367, 
        nc10368, nc10369, nc10370, nc10371, nc10372, nc10373, nc10374, 
        nc10375, nc10376, nc10377, nc10378, nc10379, 
        \B_DOUT_TEMPR88[24] , \B_DOUT_TEMPR88[23] , 
        \B_DOUT_TEMPR88[22] , \B_DOUT_TEMPR88[21] , 
        \B_DOUT_TEMPR88[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[88][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[19]  (.A(OR4_1407_Y), .B(OR4_1098_Y), .C(OR4_967_Y)
        , .D(OR4_57_Y), .Y(A_DOUT[19]));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[13]  (.A(CFG3_6_Y), .B(
        CFG3_15_Y), .Y(\BLKY2[13] ));
    OR4 OR4_537 (.A(\A_DOUT_TEMPR12[4] ), .B(\A_DOUT_TEMPR13[4] ), .C(
        \A_DOUT_TEMPR14[4] ), .D(\A_DOUT_TEMPR15[4] ), .Y(OR4_537_Y));
    OR4 OR4_1540 (.A(\A_DOUT_TEMPR32[20] ), .B(\A_DOUT_TEMPR33[20] ), 
        .C(\A_DOUT_TEMPR34[20] ), .D(\A_DOUT_TEMPR35[20] ), .Y(
        OR4_1540_Y));
    OR4 OR4_2659 (.A(\B_DOUT_TEMPR79[22] ), .B(\B_DOUT_TEMPR80[22] ), 
        .C(\B_DOUT_TEMPR81[22] ), .D(\B_DOUT_TEMPR82[22] ), .Y(
        OR4_2659_Y));
    OR4 OR4_2569 (.A(\A_DOUT_TEMPR115[10] ), .B(\A_DOUT_TEMPR116[10] ), 
        .C(\A_DOUT_TEMPR117[10] ), .D(\A_DOUT_TEMPR118[10] ), .Y(
        OR4_2569_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%46%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R46C3 (
        .A_DOUT({nc10380, nc10381, nc10382, nc10383, nc10384, nc10385, 
        nc10386, nc10387, nc10388, nc10389, nc10390, nc10391, nc10392, 
        nc10393, nc10394, \A_DOUT_TEMPR46[19] , \A_DOUT_TEMPR46[18] , 
        \A_DOUT_TEMPR46[17] , \A_DOUT_TEMPR46[16] , 
        \A_DOUT_TEMPR46[15] }), .B_DOUT({nc10395, nc10396, nc10397, 
        nc10398, nc10399, nc10400, nc10401, nc10402, nc10403, nc10404, 
        nc10405, nc10406, nc10407, nc10408, nc10409, 
        \B_DOUT_TEMPR46[19] , \B_DOUT_TEMPR46[18] , 
        \B_DOUT_TEMPR46[17] , \B_DOUT_TEMPR46[16] , 
        \B_DOUT_TEMPR46[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[46][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%32%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R32C4 (
        .A_DOUT({nc10410, nc10411, nc10412, nc10413, nc10414, nc10415, 
        nc10416, nc10417, nc10418, nc10419, nc10420, nc10421, nc10422, 
        nc10423, nc10424, \A_DOUT_TEMPR32[24] , \A_DOUT_TEMPR32[23] , 
        \A_DOUT_TEMPR32[22] , \A_DOUT_TEMPR32[21] , 
        \A_DOUT_TEMPR32[20] }), .B_DOUT({nc10425, nc10426, nc10427, 
        nc10428, nc10429, nc10430, nc10431, nc10432, nc10433, nc10434, 
        nc10435, nc10436, nc10437, nc10438, nc10439, 
        \B_DOUT_TEMPR32[24] , \B_DOUT_TEMPR32[23] , 
        \B_DOUT_TEMPR32[22] , \B_DOUT_TEMPR32[21] , 
        \B_DOUT_TEMPR32[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[32][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1159 (.A(OR4_2074_Y), .B(OR4_2368_Y), .C(OR4_2013_Y), .D(
        OR4_2386_Y), .Y(OR4_1159_Y));
    OR4 \OR4_B_DOUT[5]  (.A(OR4_811_Y), .B(OR4_1512_Y), .C(OR4_1284_Y), 
        .D(OR4_557_Y), .Y(B_DOUT[5]));
    OR4 OR4_1791 (.A(\B_DOUT_TEMPR79[25] ), .B(\B_DOUT_TEMPR80[25] ), 
        .C(\B_DOUT_TEMPR81[25] ), .D(\B_DOUT_TEMPR82[25] ), .Y(
        OR4_1791_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%2%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R2C3 (
        .A_DOUT({nc10440, nc10441, nc10442, nc10443, nc10444, nc10445, 
        nc10446, nc10447, nc10448, nc10449, nc10450, nc10451, nc10452, 
        nc10453, nc10454, \A_DOUT_TEMPR2[19] , \A_DOUT_TEMPR2[18] , 
        \A_DOUT_TEMPR2[17] , \A_DOUT_TEMPR2[16] , \A_DOUT_TEMPR2[15] })
        , .B_DOUT({nc10455, nc10456, nc10457, nc10458, nc10459, 
        nc10460, nc10461, nc10462, nc10463, nc10464, nc10465, nc10466, 
        nc10467, nc10468, nc10469, \B_DOUT_TEMPR2[19] , 
        \B_DOUT_TEMPR2[18] , \B_DOUT_TEMPR2[17] , \B_DOUT_TEMPR2[16] , 
        \B_DOUT_TEMPR2[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%1%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R1C3 (
        .A_DOUT({nc10470, nc10471, nc10472, nc10473, nc10474, nc10475, 
        nc10476, nc10477, nc10478, nc10479, nc10480, nc10481, nc10482, 
        nc10483, nc10484, \A_DOUT_TEMPR1[19] , \A_DOUT_TEMPR1[18] , 
        \A_DOUT_TEMPR1[17] , \A_DOUT_TEMPR1[16] , \A_DOUT_TEMPR1[15] })
        , .B_DOUT({nc10485, nc10486, nc10487, nc10488, nc10489, 
        nc10490, nc10491, nc10492, nc10493, nc10494, nc10495, nc10496, 
        nc10497, nc10498, nc10499, \B_DOUT_TEMPR1[19] , 
        \B_DOUT_TEMPR1[18] , \B_DOUT_TEMPR1[17] , \B_DOUT_TEMPR1[16] , 
        \B_DOUT_TEMPR1[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%96%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R96C5 (
        .A_DOUT({nc10500, nc10501, nc10502, nc10503, nc10504, nc10505, 
        nc10506, nc10507, nc10508, nc10509, nc10510, nc10511, nc10512, 
        nc10513, nc10514, \A_DOUT_TEMPR96[29] , \A_DOUT_TEMPR96[28] , 
        \A_DOUT_TEMPR96[27] , \A_DOUT_TEMPR96[26] , 
        \A_DOUT_TEMPR96[25] }), .B_DOUT({nc10515, nc10516, nc10517, 
        nc10518, nc10519, nc10520, nc10521, nc10522, nc10523, nc10524, 
        nc10525, nc10526, nc10527, nc10528, nc10529, 
        \B_DOUT_TEMPR96[29] , \B_DOUT_TEMPR96[28] , 
        \B_DOUT_TEMPR96[27] , \B_DOUT_TEMPR96[26] , 
        \B_DOUT_TEMPR96[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[96][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%99%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R99C5 (
        .A_DOUT({nc10530, nc10531, nc10532, nc10533, nc10534, nc10535, 
        nc10536, nc10537, nc10538, nc10539, nc10540, nc10541, nc10542, 
        nc10543, nc10544, \A_DOUT_TEMPR99[29] , \A_DOUT_TEMPR99[28] , 
        \A_DOUT_TEMPR99[27] , \A_DOUT_TEMPR99[26] , 
        \A_DOUT_TEMPR99[25] }), .B_DOUT({nc10545, nc10546, nc10547, 
        nc10548, nc10549, nc10550, nc10551, nc10552, nc10553, nc10554, 
        nc10555, nc10556, nc10557, nc10558, nc10559, 
        \B_DOUT_TEMPR99[29] , \B_DOUT_TEMPR99[28] , 
        \B_DOUT_TEMPR99[27] , \B_DOUT_TEMPR99[26] , 
        \B_DOUT_TEMPR99[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[99][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2534 (.A(\B_DOUT_TEMPR75[34] ), .B(\B_DOUT_TEMPR76[34] ), 
        .C(\B_DOUT_TEMPR77[34] ), .D(\B_DOUT_TEMPR78[34] ), .Y(
        OR4_2534_Y));
    OR4 OR4_1388 (.A(OR4_1557_Y), .B(OR4_499_Y), .C(OR4_2141_Y), .D(
        OR4_96_Y), .Y(OR4_1388_Y));
    OR4 OR4_2616 (.A(OR4_1153_Y), .B(OR4_2561_Y), .C(OR4_2057_Y), .D(
        OR4_1437_Y), .Y(OR4_2616_Y));
    OR4 OR4_2187 (.A(OR4_315_Y), .B(OR4_2178_Y), .C(OR4_2922_Y), .D(
        OR4_139_Y), .Y(OR4_2187_Y));
    OR4 OR4_1978 (.A(OR4_2168_Y), .B(OR4_815_Y), .C(OR4_179_Y), .D(
        OR4_2554_Y), .Y(OR4_1978_Y));
    OR4 OR4_2362 (.A(\A_DOUT_TEMPR24[24] ), .B(\A_DOUT_TEMPR25[24] ), 
        .C(\A_DOUT_TEMPR26[24] ), .D(\A_DOUT_TEMPR27[24] ), .Y(
        OR4_2362_Y));
    OR4 OR4_2110 (.A(\B_DOUT_TEMPR8[10] ), .B(\B_DOUT_TEMPR9[10] ), .C(
        \B_DOUT_TEMPR10[10] ), .D(\B_DOUT_TEMPR11[10] ), .Y(OR4_2110_Y)
        );
    OR4 OR4_2684 (.A(\A_DOUT_TEMPR48[28] ), .B(\A_DOUT_TEMPR49[28] ), 
        .C(\A_DOUT_TEMPR50[28] ), .D(\A_DOUT_TEMPR51[28] ), .Y(
        OR4_2684_Y));
    OR4 OR4_1534 (.A(\A_DOUT_TEMPR12[33] ), .B(\A_DOUT_TEMPR13[33] ), 
        .C(\A_DOUT_TEMPR14[33] ), .D(\A_DOUT_TEMPR15[33] ), .Y(
        OR4_1534_Y));
    OR4 OR4_2608 (.A(\B_DOUT_TEMPR4[0] ), .B(\B_DOUT_TEMPR5[0] ), .C(
        \B_DOUT_TEMPR6[0] ), .D(\B_DOUT_TEMPR7[0] ), .Y(OR4_2608_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%17%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R17C2 (
        .A_DOUT({nc10560, nc10561, nc10562, nc10563, nc10564, nc10565, 
        nc10566, nc10567, nc10568, nc10569, nc10570, nc10571, nc10572, 
        nc10573, nc10574, \A_DOUT_TEMPR17[14] , \A_DOUT_TEMPR17[13] , 
        \A_DOUT_TEMPR17[12] , \A_DOUT_TEMPR17[11] , 
        \A_DOUT_TEMPR17[10] }), .B_DOUT({nc10575, nc10576, nc10577, 
        nc10578, nc10579, nc10580, nc10581, nc10582, nc10583, nc10584, 
        nc10585, nc10586, nc10587, nc10588, nc10589, 
        \B_DOUT_TEMPR17[14] , \B_DOUT_TEMPR17[13] , 
        \B_DOUT_TEMPR17[12] , \B_DOUT_TEMPR17[11] , 
        \B_DOUT_TEMPR17[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_573 (.A(OR4_1567_Y), .B(OR4_2476_Y), .C(OR4_2125_Y), .D(
        OR4_589_Y), .Y(OR4_573_Y));
    OR4 OR4_286 (.A(\A_DOUT_TEMPR16[14] ), .B(\A_DOUT_TEMPR17[14] ), 
        .C(\A_DOUT_TEMPR18[14] ), .D(\A_DOUT_TEMPR19[14] ), .Y(
        OR4_286_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%113%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R113C6 (
        .A_DOUT({nc10590, nc10591, nc10592, nc10593, nc10594, nc10595, 
        nc10596, nc10597, nc10598, nc10599, nc10600, nc10601, nc10602, 
        nc10603, nc10604, \A_DOUT_TEMPR113[34] , \A_DOUT_TEMPR113[33] , 
        \A_DOUT_TEMPR113[32] , \A_DOUT_TEMPR113[31] , 
        \A_DOUT_TEMPR113[30] }), .B_DOUT({nc10605, nc10606, nc10607, 
        nc10608, nc10609, nc10610, nc10611, nc10612, nc10613, nc10614, 
        nc10615, nc10616, nc10617, nc10618, nc10619, 
        \B_DOUT_TEMPR113[34] , \B_DOUT_TEMPR113[33] , 
        \B_DOUT_TEMPR113[32] , \B_DOUT_TEMPR113[31] , 
        \B_DOUT_TEMPR113[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[113][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_294 (.A(\A_DOUT_TEMPR115[0] ), .B(\A_DOUT_TEMPR116[0] ), 
        .C(\A_DOUT_TEMPR117[0] ), .D(\A_DOUT_TEMPR118[0] ), .Y(
        OR4_294_Y));
    OR4 OR4_2240 (.A(OR4_926_Y), .B(OR4_1922_Y), .C(OR4_357_Y), .D(
        OR4_1924_Y), .Y(OR4_2240_Y));
    OR4 OR4_106 (.A(\B_DOUT_TEMPR99[0] ), .B(\B_DOUT_TEMPR100[0] ), .C(
        \B_DOUT_TEMPR101[0] ), .D(\B_DOUT_TEMPR102[0] ), .Y(OR4_106_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%59%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R59C3 (
        .A_DOUT({nc10620, nc10621, nc10622, nc10623, nc10624, nc10625, 
        nc10626, nc10627, nc10628, nc10629, nc10630, nc10631, nc10632, 
        nc10633, nc10634, \A_DOUT_TEMPR59[19] , \A_DOUT_TEMPR59[18] , 
        \A_DOUT_TEMPR59[17] , \A_DOUT_TEMPR59[16] , 
        \A_DOUT_TEMPR59[15] }), .B_DOUT({nc10635, nc10636, nc10637, 
        nc10638, nc10639, nc10640, nc10641, nc10642, nc10643, nc10644, 
        nc10645, nc10646, nc10647, nc10648, nc10649, 
        \B_DOUT_TEMPR59[19] , \B_DOUT_TEMPR59[18] , 
        \B_DOUT_TEMPR59[17] , \B_DOUT_TEMPR59[16] , 
        \B_DOUT_TEMPR59[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[59][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_412 (.A(\A_DOUT_TEMPR36[14] ), .B(\A_DOUT_TEMPR37[14] ), 
        .C(\A_DOUT_TEMPR38[14] ), .D(\A_DOUT_TEMPR39[14] ), .Y(
        OR4_412_Y));
    OR4 OR4_1945 (.A(\B_DOUT_TEMPR40[19] ), .B(\B_DOUT_TEMPR41[19] ), 
        .C(\B_DOUT_TEMPR42[19] ), .D(\B_DOUT_TEMPR43[19] ), .Y(
        OR4_1945_Y));
    OR4 OR4_790 (.A(\A_DOUT_TEMPR0[29] ), .B(\A_DOUT_TEMPR1[29] ), .C(
        \A_DOUT_TEMPR2[29] ), .D(\A_DOUT_TEMPR3[29] ), .Y(OR4_790_Y));
    OR4 OR4_1017 (.A(\B_DOUT_TEMPR68[8] ), .B(\B_DOUT_TEMPR69[8] ), .C(
        \B_DOUT_TEMPR70[8] ), .D(\B_DOUT_TEMPR71[8] ), .Y(OR4_1017_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%71%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R71C5 (
        .A_DOUT({nc10650, nc10651, nc10652, nc10653, nc10654, nc10655, 
        nc10656, nc10657, nc10658, nc10659, nc10660, nc10661, nc10662, 
        nc10663, nc10664, \A_DOUT_TEMPR71[29] , \A_DOUT_TEMPR71[28] , 
        \A_DOUT_TEMPR71[27] , \A_DOUT_TEMPR71[26] , 
        \A_DOUT_TEMPR71[25] }), .B_DOUT({nc10665, nc10666, nc10667, 
        nc10668, nc10669, nc10670, nc10671, nc10672, nc10673, nc10674, 
        nc10675, nc10676, nc10677, nc10678, nc10679, 
        \B_DOUT_TEMPR71[29] , \B_DOUT_TEMPR71[28] , 
        \B_DOUT_TEMPR71[27] , \B_DOUT_TEMPR71[26] , 
        \B_DOUT_TEMPR71[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[71][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2231 (.A(\B_DOUT_TEMPR8[36] ), .B(\B_DOUT_TEMPR9[36] ), .C(
        \B_DOUT_TEMPR10[36] ), .D(\B_DOUT_TEMPR11[36] ), .Y(OR4_2231_Y)
        );
    OR4 OR4_1319 (.A(\A_DOUT_TEMPR115[27] ), .B(\A_DOUT_TEMPR116[27] ), 
        .C(\A_DOUT_TEMPR117[27] ), .D(\A_DOUT_TEMPR118[27] ), .Y(
        OR4_1319_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%7%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R7C3 (
        .A_DOUT({nc10680, nc10681, nc10682, nc10683, nc10684, nc10685, 
        nc10686, nc10687, nc10688, nc10689, nc10690, nc10691, nc10692, 
        nc10693, nc10694, \A_DOUT_TEMPR7[19] , \A_DOUT_TEMPR7[18] , 
        \A_DOUT_TEMPR7[17] , \A_DOUT_TEMPR7[16] , \A_DOUT_TEMPR7[15] })
        , .B_DOUT({nc10695, nc10696, nc10697, nc10698, nc10699, 
        nc10700, nc10701, nc10702, nc10703, nc10704, nc10705, nc10706, 
        nc10707, nc10708, nc10709, \B_DOUT_TEMPR7[19] , 
        \B_DOUT_TEMPR7[18] , \B_DOUT_TEMPR7[17] , \B_DOUT_TEMPR7[16] , 
        \B_DOUT_TEMPR7[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1493 (.A(\A_DOUT_TEMPR4[35] ), .B(\A_DOUT_TEMPR5[35] ), .C(
        \A_DOUT_TEMPR6[35] ), .D(\A_DOUT_TEMPR7[35] ), .Y(OR4_1493_Y));
    OR4 OR4_1217 (.A(\A_DOUT_TEMPR16[3] ), .B(\A_DOUT_TEMPR17[3] ), .C(
        \A_DOUT_TEMPR18[3] ), .D(\A_DOUT_TEMPR19[3] ), .Y(OR4_1217_Y));
    OR4 OR4_2565 (.A(OR4_2291_Y), .B(OR4_1683_Y), .C(OR4_2377_Y), .D(
        OR4_2701_Y), .Y(OR4_2565_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%84%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R84C7 (
        .A_DOUT({nc10710, nc10711, nc10712, nc10713, nc10714, nc10715, 
        nc10716, nc10717, nc10718, nc10719, nc10720, nc10721, nc10722, 
        nc10723, nc10724, \A_DOUT_TEMPR84[39] , \A_DOUT_TEMPR84[38] , 
        \A_DOUT_TEMPR84[37] , \A_DOUT_TEMPR84[36] , 
        \A_DOUT_TEMPR84[35] }), .B_DOUT({nc10725, nc10726, nc10727, 
        nc10728, nc10729, nc10730, nc10731, nc10732, nc10733, nc10734, 
        nc10735, nc10736, nc10737, nc10738, nc10739, 
        \B_DOUT_TEMPR84[39] , \B_DOUT_TEMPR84[38] , 
        \B_DOUT_TEMPR84[37] , \B_DOUT_TEMPR84[36] , 
        \B_DOUT_TEMPR84[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[84][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1649 (.A(OR4_118_Y), .B(OR4_2165_Y), .C(OR4_2380_Y), .D(
        OR4_2175_Y), .Y(OR4_1649_Y));
    OR4 OR4_1231 (.A(OR4_1129_Y), .B(OR4_128_Y), .C(OR4_330_Y), .D(
        OR4_134_Y), .Y(OR4_1231_Y));
    OR4 OR4_2328 (.A(\A_DOUT_TEMPR44[1] ), .B(\A_DOUT_TEMPR45[1] ), .C(
        \A_DOUT_TEMPR46[1] ), .D(\A_DOUT_TEMPR47[1] ), .Y(OR4_2328_Y));
    OR4 OR4_1177 (.A(\A_DOUT_TEMPR60[7] ), .B(\A_DOUT_TEMPR61[7] ), .C(
        \A_DOUT_TEMPR62[7] ), .D(\A_DOUT_TEMPR63[7] ), .Y(OR4_1177_Y));
    OR4 OR4_1674 (.A(\A_DOUT_TEMPR68[35] ), .B(\A_DOUT_TEMPR69[35] ), 
        .C(\A_DOUT_TEMPR70[35] ), .D(\A_DOUT_TEMPR71[35] ), .Y(
        OR4_1674_Y));
    OR4 OR4_2346 (.A(\B_DOUT_TEMPR0[38] ), .B(\B_DOUT_TEMPR1[38] ), .C(
        \B_DOUT_TEMPR2[38] ), .D(\B_DOUT_TEMPR3[38] ), .Y(OR4_2346_Y));
    OR4 OR4_1910 (.A(\A_DOUT_TEMPR99[5] ), .B(\A_DOUT_TEMPR100[5] ), 
        .C(\A_DOUT_TEMPR101[5] ), .D(\A_DOUT_TEMPR102[5] ), .Y(
        OR4_1910_Y));
    OR4 OR4_966 (.A(\B_DOUT_TEMPR40[12] ), .B(\B_DOUT_TEMPR41[12] ), 
        .C(\B_DOUT_TEMPR42[12] ), .D(\B_DOUT_TEMPR43[12] ), .Y(
        OR4_966_Y));
    OR4 OR4_1485 (.A(\A_DOUT_TEMPR99[14] ), .B(\A_DOUT_TEMPR100[14] ), 
        .C(\A_DOUT_TEMPR101[14] ), .D(\A_DOUT_TEMPR102[14] ), .Y(
        OR4_1485_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%57%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R57C3 (
        .A_DOUT({nc10740, nc10741, nc10742, nc10743, nc10744, nc10745, 
        nc10746, nc10747, nc10748, nc10749, nc10750, nc10751, nc10752, 
        nc10753, nc10754, \A_DOUT_TEMPR57[19] , \A_DOUT_TEMPR57[18] , 
        \A_DOUT_TEMPR57[17] , \A_DOUT_TEMPR57[16] , 
        \A_DOUT_TEMPR57[15] }), .B_DOUT({nc10755, nc10756, nc10757, 
        nc10758, nc10759, nc10760, nc10761, nc10762, nc10763, nc10764, 
        nc10765, nc10766, nc10767, nc10768, nc10769, 
        \B_DOUT_TEMPR57[19] , \B_DOUT_TEMPR57[18] , 
        \B_DOUT_TEMPR57[17] , \B_DOUT_TEMPR57[16] , 
        \B_DOUT_TEMPR57[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[57][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2872 (.A(OR4_1382_Y), .B(OR4_2988_Y), .C(OR4_1142_Y), .D(
        OR4_859_Y), .Y(OR4_2872_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%64%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R64C0 (
        .A_DOUT({nc10770, nc10771, nc10772, nc10773, nc10774, nc10775, 
        nc10776, nc10777, nc10778, nc10779, nc10780, nc10781, nc10782, 
        nc10783, nc10784, \A_DOUT_TEMPR64[4] , \A_DOUT_TEMPR64[3] , 
        \A_DOUT_TEMPR64[2] , \A_DOUT_TEMPR64[1] , \A_DOUT_TEMPR64[0] })
        , .B_DOUT({nc10785, nc10786, nc10787, nc10788, nc10789, 
        nc10790, nc10791, nc10792, nc10793, nc10794, nc10795, nc10796, 
        nc10797, nc10798, nc10799, \B_DOUT_TEMPR64[4] , 
        \B_DOUT_TEMPR64[3] , \B_DOUT_TEMPR64[2] , \B_DOUT_TEMPR64[1] , 
        \B_DOUT_TEMPR64[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[64][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[33]  (.A(OR4_2182_Y), .B(OR4_1926_Y), .C(
        OR4_1035_Y), .D(OR4_1611_Y), .Y(B_DOUT[33]));
    OR4 OR4_503 (.A(\A_DOUT_TEMPR107[3] ), .B(\A_DOUT_TEMPR108[3] ), 
        .C(\A_DOUT_TEMPR109[3] ), .D(\A_DOUT_TEMPR110[3] ), .Y(
        OR4_503_Y));
    OR4 OR4_736 (.A(\A_DOUT_TEMPR87[25] ), .B(\A_DOUT_TEMPR88[25] ), 
        .C(\A_DOUT_TEMPR89[25] ), .D(\A_DOUT_TEMPR90[25] ), .Y(
        OR4_736_Y));
    OR4 OR4_2057 (.A(\A_DOUT_TEMPR111[9] ), .B(\A_DOUT_TEMPR112[9] ), 
        .C(\A_DOUT_TEMPR113[9] ), .D(\A_DOUT_TEMPR114[9] ), .Y(
        OR4_2057_Y));
    OR4 OR4_729 (.A(\A_DOUT_TEMPR91[22] ), .B(\A_DOUT_TEMPR92[22] ), 
        .C(\A_DOUT_TEMPR93[22] ), .D(\A_DOUT_TEMPR94[22] ), .Y(
        OR4_729_Y));
    OR4 OR4_12 (.A(\B_DOUT_TEMPR40[6] ), .B(\B_DOUT_TEMPR41[6] ), .C(
        \B_DOUT_TEMPR42[6] ), .D(\B_DOUT_TEMPR43[6] ), .Y(OR4_12_Y));
    OR4 OR4_2359 (.A(\B_DOUT_TEMPR68[38] ), .B(\B_DOUT_TEMPR69[38] ), 
        .C(\B_DOUT_TEMPR70[38] ), .D(\B_DOUT_TEMPR71[38] ), .Y(
        OR4_2359_Y));
    OR4 OR4_2690 (.A(OR4_2244_Y), .B(OR4_2431_Y), .C(OR4_1362_Y), .D(
        OR4_992_Y), .Y(OR4_2690_Y));
    OR4 OR4_2257 (.A(\B_DOUT_TEMPR60[16] ), .B(\B_DOUT_TEMPR61[16] ), 
        .C(\B_DOUT_TEMPR62[16] ), .D(\B_DOUT_TEMPR63[16] ), .Y(
        OR4_2257_Y));
    OR4 OR4_2098 (.A(\B_DOUT_TEMPR99[38] ), .B(\B_DOUT_TEMPR100[38] ), 
        .C(\B_DOUT_TEMPR101[38] ), .D(\B_DOUT_TEMPR102[38] ), .Y(
        OR4_2098_Y));
    OR4 OR4_1852 (.A(\A_DOUT_TEMPR52[34] ), .B(\A_DOUT_TEMPR53[34] ), 
        .C(\A_DOUT_TEMPR54[34] ), .D(\A_DOUT_TEMPR55[34] ), .Y(
        OR4_1852_Y));
    OR4 OR4_625 (.A(\A_DOUT_TEMPR115[2] ), .B(\A_DOUT_TEMPR116[2] ), 
        .C(\A_DOUT_TEMPR117[2] ), .D(\A_DOUT_TEMPR118[2] ), .Y(
        OR4_625_Y));
    OR4 OR4_1712 (.A(OR4_725_Y), .B(OR4_2818_Y), .C(OR4_3019_Y), .D(
        OR4_2834_Y), .Y(OR4_1712_Y));
    OR4 \OR4_A_DOUT[8]  (.A(OR4_388_Y), .B(OR4_2345_Y), .C(OR4_783_Y), 
        .D(OR4_281_Y), .Y(A_DOUT[8]));
    OR4 OR4_1921 (.A(\B_DOUT_TEMPR83[15] ), .B(\B_DOUT_TEMPR84[15] ), 
        .C(\B_DOUT_TEMPR85[15] ), .D(\B_DOUT_TEMPR86[15] ), .Y(
        OR4_1921_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%66%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R66C7 (
        .A_DOUT({nc10800, nc10801, nc10802, nc10803, nc10804, nc10805, 
        nc10806, nc10807, nc10808, nc10809, nc10810, nc10811, nc10812, 
        nc10813, nc10814, \A_DOUT_TEMPR66[39] , \A_DOUT_TEMPR66[38] , 
        \A_DOUT_TEMPR66[37] , \A_DOUT_TEMPR66[36] , 
        \A_DOUT_TEMPR66[35] }), .B_DOUT({nc10815, nc10816, nc10817, 
        nc10818, nc10819, nc10820, nc10821, nc10822, nc10823, nc10824, 
        nc10825, nc10826, nc10827, nc10828, nc10829, 
        \B_DOUT_TEMPR66[39] , \B_DOUT_TEMPR66[38] , 
        \B_DOUT_TEMPR66[37] , \B_DOUT_TEMPR66[36] , 
        \B_DOUT_TEMPR66[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[66][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2968 (.A(\A_DOUT_TEMPR4[11] ), .B(\A_DOUT_TEMPR5[11] ), .C(
        \A_DOUT_TEMPR6[11] ), .D(\A_DOUT_TEMPR7[11] ), .Y(OR4_2968_Y));
    OR4 OR4_989 (.A(OR4_2115_Y), .B(OR4_263_Y), .C(OR4_1331_Y), .D(
        OR4_2033_Y), .Y(OR4_989_Y));
    OR4 OR4_2913 (.A(\A_DOUT_TEMPR28[31] ), .B(\A_DOUT_TEMPR29[31] ), 
        .C(\A_DOUT_TEMPR30[31] ), .D(\A_DOUT_TEMPR31[31] ), .Y(
        OR4_2913_Y));
    OR4 OR4_1786 (.A(\A_DOUT_TEMPR52[24] ), .B(\A_DOUT_TEMPR53[24] ), 
        .C(\A_DOUT_TEMPR54[24] ), .D(\A_DOUT_TEMPR55[24] ), .Y(
        OR4_1786_Y));
    OR4 OR4_229 (.A(\A_DOUT_TEMPR4[14] ), .B(\A_DOUT_TEMPR5[14] ), .C(
        \A_DOUT_TEMPR6[14] ), .D(\A_DOUT_TEMPR7[14] ), .Y(OR4_229_Y));
    OR4 OR4_2950 (.A(OR4_79_Y), .B(OR4_1577_Y), .C(OR4_2143_Y), .D(
        OR4_1967_Y), .Y(OR4_2950_Y));
    OR4 OR4_2673 (.A(\B_DOUT_TEMPR79[4] ), .B(\B_DOUT_TEMPR80[4] ), .C(
        \B_DOUT_TEMPR81[4] ), .D(\B_DOUT_TEMPR82[4] ), .Y(OR4_2673_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%39%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R39C3 (
        .A_DOUT({nc10830, nc10831, nc10832, nc10833, nc10834, nc10835, 
        nc10836, nc10837, nc10838, nc10839, nc10840, nc10841, nc10842, 
        nc10843, nc10844, \A_DOUT_TEMPR39[19] , \A_DOUT_TEMPR39[18] , 
        \A_DOUT_TEMPR39[17] , \A_DOUT_TEMPR39[16] , 
        \A_DOUT_TEMPR39[15] }), .B_DOUT({nc10845, nc10846, nc10847, 
        nc10848, nc10849, nc10850, nc10851, nc10852, nc10853, nc10854, 
        nc10855, nc10856, nc10857, nc10858, nc10859, 
        \B_DOUT_TEMPR39[19] , \B_DOUT_TEMPR39[18] , 
        \B_DOUT_TEMPR39[17] , \B_DOUT_TEMPR39[16] , 
        \B_DOUT_TEMPR39[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[39][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%67%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R67C6 (
        .A_DOUT({nc10860, nc10861, nc10862, nc10863, nc10864, nc10865, 
        nc10866, nc10867, nc10868, nc10869, nc10870, nc10871, nc10872, 
        nc10873, nc10874, \A_DOUT_TEMPR67[34] , \A_DOUT_TEMPR67[33] , 
        \A_DOUT_TEMPR67[32] , \A_DOUT_TEMPR67[31] , 
        \A_DOUT_TEMPR67[30] }), .B_DOUT({nc10875, nc10876, nc10877, 
        nc10878, nc10879, nc10880, nc10881, nc10882, nc10883, nc10884, 
        nc10885, nc10886, nc10887, nc10888, nc10889, 
        \B_DOUT_TEMPR67[34] , \B_DOUT_TEMPR67[33] , 
        \B_DOUT_TEMPR67[32] , \B_DOUT_TEMPR67[31] , 
        \B_DOUT_TEMPR67[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[67][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2979 (.A(OR4_1982_Y), .B(OR4_2357_Y), .C(OR4_73_Y), .D(
        OR4_904_Y), .Y(OR4_2979_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%2%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R2C7 (
        .A_DOUT({nc10890, nc10891, nc10892, nc10893, nc10894, nc10895, 
        nc10896, nc10897, nc10898, nc10899, nc10900, nc10901, nc10902, 
        nc10903, nc10904, \A_DOUT_TEMPR2[39] , \A_DOUT_TEMPR2[38] , 
        \A_DOUT_TEMPR2[37] , \A_DOUT_TEMPR2[36] , \A_DOUT_TEMPR2[35] })
        , .B_DOUT({nc10905, nc10906, nc10907, nc10908, nc10909, 
        nc10910, nc10911, nc10912, nc10913, nc10914, nc10915, nc10916, 
        nc10917, nc10918, nc10919, \B_DOUT_TEMPR2[39] , 
        \B_DOUT_TEMPR2[38] , \B_DOUT_TEMPR2[37] , \B_DOUT_TEMPR2[36] , 
        \B_DOUT_TEMPR2[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_723 (.A(OR4_955_Y), .B(OR4_2111_Y), .C(OR2_3_Y), .D(
        \B_DOUT_TEMPR74[17] ), .Y(OR4_723_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENB[2]  (.A(B_WBYTE_EN[1]), .B(
        B_WEN), .Y(\WBYTEENB[2] ));
    OR4 OR4_2425 (.A(\A_DOUT_TEMPR12[15] ), .B(\A_DOUT_TEMPR13[15] ), 
        .C(\A_DOUT_TEMPR14[15] ), .D(\A_DOUT_TEMPR15[15] ), .Y(
        OR4_2425_Y));
    OR4 OR4_531 (.A(\A_DOUT_TEMPR20[28] ), .B(\A_DOUT_TEMPR21[28] ), 
        .C(\A_DOUT_TEMPR22[28] ), .D(\A_DOUT_TEMPR23[28] ), .Y(
        OR4_531_Y));
    OR4 OR4_2680 (.A(\B_DOUT_TEMPR87[37] ), .B(\B_DOUT_TEMPR88[37] ), 
        .C(\B_DOUT_TEMPR89[37] ), .D(\B_DOUT_TEMPR90[37] ), .Y(
        OR4_2680_Y));
    OR4 OR4_538 (.A(\A_DOUT_TEMPR16[20] ), .B(\A_DOUT_TEMPR17[20] ), 
        .C(\A_DOUT_TEMPR18[20] ), .D(\A_DOUT_TEMPR19[20] ), .Y(
        OR4_538_Y));
    OR4 OR4_1004 (.A(\A_DOUT_TEMPR68[37] ), .B(\A_DOUT_TEMPR69[37] ), 
        .C(\A_DOUT_TEMPR70[37] ), .D(\A_DOUT_TEMPR71[37] ), .Y(
        OR4_1004_Y));
    OR4 OR4_1006 (.A(\A_DOUT_TEMPR60[21] ), .B(\A_DOUT_TEMPR61[21] ), 
        .C(\A_DOUT_TEMPR62[21] ), .D(\A_DOUT_TEMPR63[21] ), .Y(
        OR4_1006_Y));
    OR4 OR4_1612 (.A(\A_DOUT_TEMPR48[16] ), .B(\A_DOUT_TEMPR49[16] ), 
        .C(\A_DOUT_TEMPR50[16] ), .D(\A_DOUT_TEMPR51[16] ), .Y(
        OR4_1612_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%62%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R62C4 (
        .A_DOUT({nc10920, nc10921, nc10922, nc10923, nc10924, nc10925, 
        nc10926, nc10927, nc10928, nc10929, nc10930, nc10931, nc10932, 
        nc10933, nc10934, \A_DOUT_TEMPR62[24] , \A_DOUT_TEMPR62[23] , 
        \A_DOUT_TEMPR62[22] , \A_DOUT_TEMPR62[21] , 
        \A_DOUT_TEMPR62[20] }), .B_DOUT({nc10935, nc10936, nc10937, 
        nc10938, nc10939, nc10940, nc10941, nc10942, nc10943, nc10944, 
        nc10945, nc10946, nc10947, nc10948, nc10949, 
        \B_DOUT_TEMPR62[24] , \B_DOUT_TEMPR62[23] , 
        \B_DOUT_TEMPR62[22] , \B_DOUT_TEMPR62[21] , 
        \B_DOUT_TEMPR62[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[62][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[28]  (.A(OR4_2466_Y), .B(OR4_605_Y), .C(OR4_2333_Y)
        , .D(OR4_1201_Y), .Y(B_DOUT[28]));
    OR4 OR4_2311 (.A(\A_DOUT_TEMPR64[18] ), .B(\A_DOUT_TEMPR65[18] ), 
        .C(\A_DOUT_TEMPR66[18] ), .D(\A_DOUT_TEMPR67[18] ), .Y(
        OR4_2311_Y));
    OR4 OR4_2088 (.A(\B_DOUT_TEMPR87[34] ), .B(\B_DOUT_TEMPR88[34] ), 
        .C(\B_DOUT_TEMPR89[34] ), .D(\B_DOUT_TEMPR90[34] ), .Y(
        OR4_2088_Y));
    OR4 OR4_2809 (.A(OR4_2612_Y), .B(OR4_2751_Y), .C(OR4_309_Y), .D(
        OR4_2546_Y), .Y(OR4_2809_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%40%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R40C0 (
        .A_DOUT({nc10950, nc10951, nc10952, nc10953, nc10954, nc10955, 
        nc10956, nc10957, nc10958, nc10959, nc10960, nc10961, nc10962, 
        nc10963, nc10964, \A_DOUT_TEMPR40[4] , \A_DOUT_TEMPR40[3] , 
        \A_DOUT_TEMPR40[2] , \A_DOUT_TEMPR40[1] , \A_DOUT_TEMPR40[0] })
        , .B_DOUT({nc10965, nc10966, nc10967, nc10968, nc10969, 
        nc10970, nc10971, nc10972, nc10973, nc10974, nc10975, nc10976, 
        nc10977, nc10978, nc10979, \B_DOUT_TEMPR40[4] , 
        \B_DOUT_TEMPR40[3] , \B_DOUT_TEMPR40[2] , \B_DOUT_TEMPR40[1] , 
        \B_DOUT_TEMPR40[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[40][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_38 (.A(OR4_2541_Y), .B(OR4_1731_Y), .C(OR4_2367_Y), .D(
        OR4_1565_Y), .Y(OR4_38_Y));
    OR4 OR4_1653 (.A(\A_DOUT_TEMPR44[30] ), .B(\A_DOUT_TEMPR45[30] ), 
        .C(\A_DOUT_TEMPR46[30] ), .D(\A_DOUT_TEMPR47[30] ), .Y(
        OR4_1653_Y));
    OR4 OR4_2442 (.A(\B_DOUT_TEMPR28[12] ), .B(\B_DOUT_TEMPR29[12] ), 
        .C(\B_DOUT_TEMPR30[12] ), .D(\B_DOUT_TEMPR31[12] ), .Y(
        OR4_2442_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%45%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R45C4 (
        .A_DOUT({nc10980, nc10981, nc10982, nc10983, nc10984, nc10985, 
        nc10986, nc10987, nc10988, nc10989, nc10990, nc10991, nc10992, 
        nc10993, nc10994, \A_DOUT_TEMPR45[24] , \A_DOUT_TEMPR45[23] , 
        \A_DOUT_TEMPR45[22] , \A_DOUT_TEMPR45[21] , 
        \A_DOUT_TEMPR45[20] }), .B_DOUT({nc10995, nc10996, nc10997, 
        nc10998, nc10999, nc11000, nc11001, nc11002, nc11003, nc11004, 
        nc11005, nc11006, nc11007, nc11008, nc11009, 
        \B_DOUT_TEMPR45[24] , \B_DOUT_TEMPR45[23] , 
        \B_DOUT_TEMPR45[22] , \B_DOUT_TEMPR45[21] , 
        \B_DOUT_TEMPR45[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%6%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R6C3 (
        .A_DOUT({nc11010, nc11011, nc11012, nc11013, nc11014, nc11015, 
        nc11016, nc11017, nc11018, nc11019, nc11020, nc11021, nc11022, 
        nc11023, nc11024, \A_DOUT_TEMPR6[19] , \A_DOUT_TEMPR6[18] , 
        \A_DOUT_TEMPR6[17] , \A_DOUT_TEMPR6[16] , \A_DOUT_TEMPR6[15] })
        , .B_DOUT({nc11025, nc11026, nc11027, nc11028, nc11029, 
        nc11030, nc11031, nc11032, nc11033, nc11034, nc11035, nc11036, 
        nc11037, nc11038, nc11039, \B_DOUT_TEMPR6[19] , 
        \B_DOUT_TEMPR6[18] , \B_DOUT_TEMPR6[17] , \B_DOUT_TEMPR6[16] , 
        \B_DOUT_TEMPR6[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2752 (.A(OR4_2272_Y), .B(OR4_1513_Y), .C(OR4_1279_Y), .D(
        OR4_763_Y), .Y(OR4_2752_Y));
    OR4 OR4_2811 (.A(OR4_1884_Y), .B(OR4_820_Y), .C(OR4_2468_Y), .D(
        OR4_419_Y), .Y(OR4_2811_Y));
    OR4 OR4_156 (.A(OR4_2060_Y), .B(OR4_1525_Y), .C(OR4_2692_Y), .D(
        OR4_2870_Y), .Y(OR4_156_Y));
    OR4 OR4_228 (.A(\A_DOUT_TEMPR8[3] ), .B(\A_DOUT_TEMPR9[3] ), .C(
        \A_DOUT_TEMPR10[3] ), .D(\A_DOUT_TEMPR11[3] ), .Y(OR4_228_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%37%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R37C3 (
        .A_DOUT({nc11040, nc11041, nc11042, nc11043, nc11044, nc11045, 
        nc11046, nc11047, nc11048, nc11049, nc11050, nc11051, nc11052, 
        nc11053, nc11054, \A_DOUT_TEMPR37[19] , \A_DOUT_TEMPR37[18] , 
        \A_DOUT_TEMPR37[17] , \A_DOUT_TEMPR37[16] , 
        \A_DOUT_TEMPR37[15] }), .B_DOUT({nc11055, nc11056, nc11057, 
        nc11058, nc11059, nc11060, nc11061, nc11062, nc11063, nc11064, 
        nc11065, nc11066, nc11067, nc11068, nc11069, 
        \B_DOUT_TEMPR37[19] , \B_DOUT_TEMPR37[18] , 
        \B_DOUT_TEMPR37[17] , \B_DOUT_TEMPR37[16] , 
        \B_DOUT_TEMPR37[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[37][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1959 (.A(\A_DOUT_TEMPR16[0] ), .B(\A_DOUT_TEMPR17[0] ), .C(
        \A_DOUT_TEMPR18[0] ), .D(\A_DOUT_TEMPR19[0] ), .Y(OR4_1959_Y));
    OR4 OR4_2448 (.A(\A_DOUT_TEMPR87[14] ), .B(\A_DOUT_TEMPR88[14] ), 
        .C(\A_DOUT_TEMPR89[14] ), .D(\A_DOUT_TEMPR90[14] ), .Y(
        OR4_2448_Y));
    OR4 OR4_1912 (.A(\B_DOUT_TEMPR91[39] ), .B(\B_DOUT_TEMPR92[39] ), 
        .C(\B_DOUT_TEMPR93[39] ), .D(\B_DOUT_TEMPR94[39] ), .Y(
        OR4_1912_Y));
    OR4 OR4_1223 (.A(\A_DOUT_TEMPR115[34] ), .B(\A_DOUT_TEMPR116[34] ), 
        .C(\A_DOUT_TEMPR117[34] ), .D(\A_DOUT_TEMPR118[34] ), .Y(
        OR4_1223_Y));
    OR4 OR4_2774 (.A(OR4_2712_Y), .B(OR4_1097_Y), .C(OR2_16_Y), .D(
        \A_DOUT_TEMPR74[9] ), .Y(OR4_2774_Y));
    OR4 OR4_2167 (.A(\B_DOUT_TEMPR0[32] ), .B(\B_DOUT_TEMPR1[32] ), .C(
        \B_DOUT_TEMPR2[32] ), .D(\B_DOUT_TEMPR3[32] ), .Y(OR4_2167_Y));
    OR4 OR4_2194 (.A(\B_DOUT_TEMPR83[1] ), .B(\B_DOUT_TEMPR84[1] ), .C(
        \B_DOUT_TEMPR85[1] ), .D(\B_DOUT_TEMPR86[1] ), .Y(OR4_2194_Y));
    OR4 OR4_2101 (.A(\B_DOUT_TEMPR52[21] ), .B(\B_DOUT_TEMPR53[21] ), 
        .C(\B_DOUT_TEMPR54[21] ), .D(\B_DOUT_TEMPR55[21] ), .Y(
        OR4_2101_Y));
    OR4 OR4_1303 (.A(\A_DOUT_TEMPR12[21] ), .B(\A_DOUT_TEMPR13[21] ), 
        .C(\A_DOUT_TEMPR14[21] ), .D(\A_DOUT_TEMPR15[21] ), .Y(
        OR4_1303_Y));
    OR4 OR4_1047 (.A(\A_DOUT_TEMPR79[32] ), .B(\A_DOUT_TEMPR80[32] ), 
        .C(\A_DOUT_TEMPR81[32] ), .D(\A_DOUT_TEMPR82[32] ), .Y(
        OR4_1047_Y));
    OR4 OR4_2664 (.A(\B_DOUT_TEMPR68[11] ), .B(\B_DOUT_TEMPR69[11] ), 
        .C(\B_DOUT_TEMPR70[11] ), .D(\B_DOUT_TEMPR71[11] ), .Y(
        OR4_2664_Y));
    OR4 OR4_2471 (.A(OR4_2990_Y), .B(OR4_2564_Y), .C(OR4_142_Y), .D(
        OR4_2371_Y), .Y(OR4_2471_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%117%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R117C1 (
        .A_DOUT({nc11070, nc11071, nc11072, nc11073, nc11074, nc11075, 
        nc11076, nc11077, nc11078, nc11079, nc11080, nc11081, nc11082, 
        nc11083, nc11084, \A_DOUT_TEMPR117[9] , \A_DOUT_TEMPR117[8] , 
        \A_DOUT_TEMPR117[7] , \A_DOUT_TEMPR117[6] , 
        \A_DOUT_TEMPR117[5] }), .B_DOUT({nc11085, nc11086, nc11087, 
        nc11088, nc11089, nc11090, nc11091, nc11092, nc11093, nc11094, 
        nc11095, nc11096, nc11097, nc11098, nc11099, 
        \B_DOUT_TEMPR117[9] , \B_DOUT_TEMPR117[8] , 
        \B_DOUT_TEMPR117[7] , \B_DOUT_TEMPR117[6] , 
        \B_DOUT_TEMPR117[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[117][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%28%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R28C0 (
        .A_DOUT({nc11100, nc11101, nc11102, nc11103, nc11104, nc11105, 
        nc11106, nc11107, nc11108, nc11109, nc11110, nc11111, nc11112, 
        nc11113, nc11114, \A_DOUT_TEMPR28[4] , \A_DOUT_TEMPR28[3] , 
        \A_DOUT_TEMPR28[2] , \A_DOUT_TEMPR28[1] , \A_DOUT_TEMPR28[0] })
        , .B_DOUT({nc11115, nc11116, nc11117, nc11118, nc11119, 
        nc11120, nc11121, nc11122, nc11123, nc11124, nc11125, nc11126, 
        nc11127, nc11128, nc11129, \B_DOUT_TEMPR28[4] , 
        \B_DOUT_TEMPR28[3] , \B_DOUT_TEMPR28[2] , \B_DOUT_TEMPR28[1] , 
        \B_DOUT_TEMPR28[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_335 (.A(\B_DOUT_TEMPR52[7] ), .B(\B_DOUT_TEMPR53[7] ), .C(
        \B_DOUT_TEMPR54[7] ), .D(\B_DOUT_TEMPR55[7] ), .Y(OR4_335_Y));
    OR4 OR4_1349 (.A(\B_DOUT_TEMPR44[36] ), .B(\B_DOUT_TEMPR45[36] ), 
        .C(\B_DOUT_TEMPR46[36] ), .D(\B_DOUT_TEMPR47[36] ), .Y(
        OR4_1349_Y));
    OR4 OR4_2726 (.A(OR4_2016_Y), .B(OR4_284_Y), .C(OR4_2989_Y), .D(
        OR4_1015_Y), .Y(OR4_2726_Y));
    OR4 OR4_1247 (.A(\A_DOUT_TEMPR75[19] ), .B(\A_DOUT_TEMPR76[19] ), 
        .C(\A_DOUT_TEMPR77[19] ), .D(\A_DOUT_TEMPR78[19] ), .Y(
        OR4_1247_Y));
    OR4 OR4_749 (.A(\A_DOUT_TEMPR95[35] ), .B(\A_DOUT_TEMPR96[35] ), 
        .C(\A_DOUT_TEMPR97[35] ), .D(\A_DOUT_TEMPR98[35] ), .Y(
        OR4_749_Y));
    OR4 OR4_14 (.A(OR4_524_Y), .B(OR4_432_Y), .C(OR4_1923_Y), .D(
        OR4_435_Y), .Y(OR4_14_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENA[10]  (.A(A_WBYTE_EN[5]), .B(
        A_WEN), .Y(\WBYTEENA[10] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%56%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R56C5 (
        .A_DOUT({nc11130, nc11131, nc11132, nc11133, nc11134, nc11135, 
        nc11136, nc11137, nc11138, nc11139, nc11140, nc11141, nc11142, 
        nc11143, nc11144, \A_DOUT_TEMPR56[29] , \A_DOUT_TEMPR56[28] , 
        \A_DOUT_TEMPR56[27] , \A_DOUT_TEMPR56[26] , 
        \A_DOUT_TEMPR56[25] }), .B_DOUT({nc11145, nc11146, nc11147, 
        nc11148, nc11149, nc11150, nc11151, nc11152, nc11153, nc11154, 
        nc11155, nc11156, nc11157, nc11158, nc11159, 
        \B_DOUT_TEMPR56[29] , \B_DOUT_TEMPR56[28] , 
        \B_DOUT_TEMPR56[27] , \B_DOUT_TEMPR56[26] , 
        \B_DOUT_TEMPR56[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[56][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%59%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R59C5 (
        .A_DOUT({nc11160, nc11161, nc11162, nc11163, nc11164, nc11165, 
        nc11166, nc11167, nc11168, nc11169, nc11170, nc11171, nc11172, 
        nc11173, nc11174, \A_DOUT_TEMPR59[29] , \A_DOUT_TEMPR59[28] , 
        \A_DOUT_TEMPR59[27] , \A_DOUT_TEMPR59[26] , 
        \A_DOUT_TEMPR59[25] }), .B_DOUT({nc11175, nc11176, nc11177, 
        nc11178, nc11179, nc11180, nc11181, nc11182, nc11183, nc11184, 
        nc11185, nc11186, nc11187, nc11188, nc11189, 
        \B_DOUT_TEMPR59[29] , \B_DOUT_TEMPR59[28] , 
        \B_DOUT_TEMPR59[27] , \B_DOUT_TEMPR59[26] , 
        \B_DOUT_TEMPR59[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[59][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2005 (.A(\B_DOUT_TEMPR48[1] ), .B(\B_DOUT_TEMPR49[1] ), .C(
        \B_DOUT_TEMPR50[1] ), .D(\B_DOUT_TEMPR51[1] ), .Y(OR4_2005_Y));
    OR4 OR4_1296 (.A(\B_DOUT_TEMPR4[10] ), .B(\B_DOUT_TEMPR5[10] ), .C(
        \B_DOUT_TEMPR6[10] ), .D(\B_DOUT_TEMPR7[10] ), .Y(OR4_1296_Y));
    OR4 OR4_2652 (.A(\B_DOUT_TEMPR20[9] ), .B(\B_DOUT_TEMPR21[9] ), .C(
        \B_DOUT_TEMPR22[9] ), .D(\B_DOUT_TEMPR23[9] ), .Y(OR4_2652_Y));
    OR4 OR4_2540 (.A(\B_DOUT_TEMPR4[1] ), .B(\B_DOUT_TEMPR5[1] ), .C(
        \B_DOUT_TEMPR6[1] ), .D(\B_DOUT_TEMPR7[1] ), .Y(OR4_2540_Y));
    OR4 OR4_1670 (.A(\A_DOUT_TEMPR52[5] ), .B(\A_DOUT_TEMPR53[5] ), .C(
        \A_DOUT_TEMPR54[5] ), .D(\A_DOUT_TEMPR55[5] ), .Y(OR4_1670_Y));
    OR4 OR4_645 (.A(\B_DOUT_TEMPR64[15] ), .B(\B_DOUT_TEMPR65[15] ), 
        .C(\B_DOUT_TEMPR66[15] ), .D(\B_DOUT_TEMPR67[15] ), .Y(
        OR4_645_Y));
    OR4 OR4_1754 (.A(\A_DOUT_TEMPR91[31] ), .B(\A_DOUT_TEMPR92[31] ), 
        .C(\A_DOUT_TEMPR93[31] ), .D(\A_DOUT_TEMPR94[31] ), .Y(
        OR4_1754_Y));
    OR4 OR4_1940 (.A(\A_DOUT_TEMPR91[1] ), .B(\A_DOUT_TEMPR92[1] ), .C(
        \A_DOUT_TEMPR93[1] ), .D(\A_DOUT_TEMPR94[1] ), .Y(OR4_1940_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%114%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R114C5 (
        .A_DOUT({nc11190, nc11191, nc11192, nc11193, nc11194, nc11195, 
        nc11196, nc11197, nc11198, nc11199, nc11200, nc11201, nc11202, 
        nc11203, nc11204, \A_DOUT_TEMPR114[29] , \A_DOUT_TEMPR114[28] , 
        \A_DOUT_TEMPR114[27] , \A_DOUT_TEMPR114[26] , 
        \A_DOUT_TEMPR114[25] }), .B_DOUT({nc11205, nc11206, nc11207, 
        nc11208, nc11209, nc11210, nc11211, nc11212, nc11213, nc11214, 
        nc11215, nc11216, nc11217, nc11218, nc11219, 
        \B_DOUT_TEMPR114[29] , \B_DOUT_TEMPR114[28] , 
        \B_DOUT_TEMPR114[27] , \B_DOUT_TEMPR114[26] , 
        \B_DOUT_TEMPR114[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[114][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_462 (.A(\A_DOUT_TEMPR20[39] ), .B(\A_DOUT_TEMPR21[39] ), 
        .C(\A_DOUT_TEMPR22[39] ), .D(\A_DOUT_TEMPR23[39] ), .Y(
        OR4_462_Y));
    OR4 OR4_1451 (.A(\B_DOUT_TEMPR20[1] ), .B(\B_DOUT_TEMPR21[1] ), .C(
        \B_DOUT_TEMPR22[1] ), .D(\B_DOUT_TEMPR23[1] ), .Y(OR4_1451_Y));
    OR4 OR4_1078 (.A(\A_DOUT_TEMPR91[6] ), .B(\A_DOUT_TEMPR92[6] ), .C(
        \A_DOUT_TEMPR93[6] ), .D(\A_DOUT_TEMPR94[6] ), .Y(OR4_1078_Y));
    OR4 OR4_249 (.A(\B_DOUT_TEMPR91[30] ), .B(\B_DOUT_TEMPR92[30] ), 
        .C(\B_DOUT_TEMPR93[30] ), .D(\B_DOUT_TEMPR94[30] ), .Y(
        OR4_249_Y));
    OR4 OR4_2952 (.A(\A_DOUT_TEMPR4[32] ), .B(\A_DOUT_TEMPR5[32] ), .C(
        \A_DOUT_TEMPR6[32] ), .D(\A_DOUT_TEMPR7[32] ), .Y(OR4_2952_Y));
    OR4 OR4_22 (.A(\A_DOUT_TEMPR28[1] ), .B(\A_DOUT_TEMPR29[1] ), .C(
        \A_DOUT_TEMPR30[1] ), .D(\A_DOUT_TEMPR31[1] ), .Y(OR4_22_Y));
    OR4 OR4_553 (.A(\B_DOUT_TEMPR56[32] ), .B(\B_DOUT_TEMPR57[32] ), 
        .C(\B_DOUT_TEMPR58[32] ), .D(\B_DOUT_TEMPR59[32] ), .Y(
        OR4_553_Y));
    OR4 OR4_2184 (.A(\B_DOUT_TEMPR40[11] ), .B(\B_DOUT_TEMPR41[11] ), 
        .C(\B_DOUT_TEMPR42[11] ), .D(\B_DOUT_TEMPR43[11] ), .Y(
        OR4_2184_Y));
    OR4 OR4_127 (.A(OR4_3038_Y), .B(OR4_919_Y), .C(OR4_553_Y), .D(
        OR4_2046_Y), .Y(OR4_127_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%83%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R83C4 (
        .A_DOUT({nc11220, nc11221, nc11222, nc11223, nc11224, nc11225, 
        nc11226, nc11227, nc11228, nc11229, nc11230, nc11231, nc11232, 
        nc11233, nc11234, \A_DOUT_TEMPR83[24] , \A_DOUT_TEMPR83[23] , 
        \A_DOUT_TEMPR83[22] , \A_DOUT_TEMPR83[21] , 
        \A_DOUT_TEMPR83[20] }), .B_DOUT({nc11235, nc11236, nc11237, 
        nc11238, nc11239, nc11240, nc11241, nc11242, nc11243, nc11244, 
        nc11245, nc11246, nc11247, nc11248, nc11249, 
        \B_DOUT_TEMPR83[24] , \B_DOUT_TEMPR83[23] , 
        \B_DOUT_TEMPR83[22] , \B_DOUT_TEMPR83[21] , 
        \B_DOUT_TEMPR83[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[83][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2895 (.A(\A_DOUT_TEMPR64[30] ), .B(\A_DOUT_TEMPR65[30] ), 
        .C(\A_DOUT_TEMPR66[30] ), .D(\A_DOUT_TEMPR67[30] ), .Y(
        OR4_2895_Y));
    OR4 OR4_743 (.A(\B_DOUT_TEMPR95[7] ), .B(\B_DOUT_TEMPR96[7] ), .C(
        \B_DOUT_TEMPR97[7] ), .D(\B_DOUT_TEMPR98[7] ), .Y(OR4_743_Y));
    OR4 OR4_2807 (.A(OR4_2597_Y), .B(OR4_987_Y), .C(OR4_460_Y), .D(
        OR4_1265_Y), .Y(OR4_2807_Y));
    OR4 OR4_2974 (.A(\A_DOUT_TEMPR20[1] ), .B(\A_DOUT_TEMPR21[1] ), .C(
        \A_DOUT_TEMPR22[1] ), .D(\A_DOUT_TEMPR23[1] ), .Y(OR4_2974_Y));
    OR4 OR4_830 (.A(\A_DOUT_TEMPR12[12] ), .B(\A_DOUT_TEMPR13[12] ), 
        .C(\A_DOUT_TEMPR14[12] ), .D(\A_DOUT_TEMPR15[12] ), .Y(
        OR4_830_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%76%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R76C3 (
        .A_DOUT({nc11250, nc11251, nc11252, nc11253, nc11254, nc11255, 
        nc11256, nc11257, nc11258, nc11259, nc11260, nc11261, nc11262, 
        nc11263, nc11264, \A_DOUT_TEMPR76[19] , \A_DOUT_TEMPR76[18] , 
        \A_DOUT_TEMPR76[17] , \A_DOUT_TEMPR76[16] , 
        \A_DOUT_TEMPR76[15] }), .B_DOUT({nc11265, nc11266, nc11267, 
        nc11268, nc11269, nc11270, nc11271, nc11272, nc11273, nc11274, 
        nc11275, nc11276, nc11277, nc11278, nc11279, 
        \B_DOUT_TEMPR76[19] , \B_DOUT_TEMPR76[18] , 
        \B_DOUT_TEMPR76[17] , \B_DOUT_TEMPR76[16] , 
        \B_DOUT_TEMPR76[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[76][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1742 (.A(\A_DOUT_TEMPR36[36] ), .B(\A_DOUT_TEMPR37[36] ), 
        .C(\A_DOUT_TEMPR38[36] ), .D(\A_DOUT_TEMPR39[36] ), .Y(
        OR4_1742_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%117%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R117C0 (
        .A_DOUT({nc11280, nc11281, nc11282, nc11283, nc11284, nc11285, 
        nc11286, nc11287, nc11288, nc11289, nc11290, nc11291, nc11292, 
        nc11293, nc11294, \A_DOUT_TEMPR117[4] , \A_DOUT_TEMPR117[3] , 
        \A_DOUT_TEMPR117[2] , \A_DOUT_TEMPR117[1] , 
        \A_DOUT_TEMPR117[0] }), .B_DOUT({nc11295, nc11296, nc11297, 
        nc11298, nc11299, nc11300, nc11301, nc11302, nc11303, nc11304, 
        nc11305, nc11306, nc11307, nc11308, nc11309, 
        \B_DOUT_TEMPR117[4] , \B_DOUT_TEMPR117[3] , 
        \B_DOUT_TEMPR117[2] , \B_DOUT_TEMPR117[1] , 
        \B_DOUT_TEMPR117[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[117][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_530 (.A(\B_DOUT_TEMPR103[16] ), .B(\B_DOUT_TEMPR104[16] ), 
        .C(\B_DOUT_TEMPR105[16] ), .D(\B_DOUT_TEMPR106[16] ), .Y(
        OR4_530_Y));
    OR4 OR4_674 (.A(\A_DOUT_TEMPR36[30] ), .B(\A_DOUT_TEMPR37[30] ), 
        .C(\A_DOUT_TEMPR38[30] ), .D(\A_DOUT_TEMPR39[30] ), .Y(
        OR4_674_Y));
    OR4 OR4_1587 (.A(\B_DOUT_TEMPR83[4] ), .B(\B_DOUT_TEMPR84[4] ), .C(
        \B_DOUT_TEMPR85[4] ), .D(\B_DOUT_TEMPR86[4] ), .Y(OR4_1587_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%14%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R14C0 (
        .A_DOUT({nc11310, nc11311, nc11312, nc11313, nc11314, nc11315, 
        nc11316, nc11317, nc11318, nc11319, nc11320, nc11321, nc11322, 
        nc11323, nc11324, \A_DOUT_TEMPR14[4] , \A_DOUT_TEMPR14[3] , 
        \A_DOUT_TEMPR14[2] , \A_DOUT_TEMPR14[1] , \A_DOUT_TEMPR14[0] })
        , .B_DOUT({nc11325, nc11326, nc11327, nc11328, nc11329, 
        nc11330, nc11331, nc11332, nc11333, nc11334, nc11335, nc11336, 
        nc11337, nc11338, nc11339, \B_DOUT_TEMPR14[4] , 
        \B_DOUT_TEMPR14[3] , \B_DOUT_TEMPR14[2] , \B_DOUT_TEMPR14[1] , 
        \B_DOUT_TEMPR14[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2976 (.A(\B_DOUT_TEMPR103[36] ), .B(\B_DOUT_TEMPR104[36] ), 
        .C(\B_DOUT_TEMPR105[36] ), .D(\B_DOUT_TEMPR106[36] ), .Y(
        OR4_2976_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%25%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R25C0 (
        .A_DOUT({nc11340, nc11341, nc11342, nc11343, nc11344, nc11345, 
        nc11346, nc11347, nc11348, nc11349, nc11350, nc11351, nc11352, 
        nc11353, nc11354, \A_DOUT_TEMPR25[4] , \A_DOUT_TEMPR25[3] , 
        \A_DOUT_TEMPR25[2] , \A_DOUT_TEMPR25[1] , \A_DOUT_TEMPR25[0] })
        , .B_DOUT({nc11355, nc11356, nc11357, nc11358, nc11359, 
        nc11360, nc11361, nc11362, nc11363, nc11364, nc11365, nc11366, 
        nc11367, nc11368, nc11369, \B_DOUT_TEMPR25[4] , 
        \B_DOUT_TEMPR25[3] , \B_DOUT_TEMPR25[2] , \B_DOUT_TEMPR25[1] , 
        \B_DOUT_TEMPR25[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_88 (.A(\A_DOUT_TEMPR4[13] ), .B(\A_DOUT_TEMPR5[13] ), .C(
        \A_DOUT_TEMPR6[13] ), .D(\A_DOUT_TEMPR7[13] ), .Y(OR4_88_Y));
    OR4 OR4_248 (.A(\B_DOUT_TEMPR87[32] ), .B(\B_DOUT_TEMPR88[32] ), 
        .C(\B_DOUT_TEMPR89[32] ), .D(\B_DOUT_TEMPR90[32] ), .Y(
        OR4_248_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%104%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R104C0 (
        .A_DOUT({nc11370, nc11371, nc11372, nc11373, nc11374, nc11375, 
        nc11376, nc11377, nc11378, nc11379, nc11380, nc11381, nc11382, 
        nc11383, nc11384, \A_DOUT_TEMPR104[4] , \A_DOUT_TEMPR104[3] , 
        \A_DOUT_TEMPR104[2] , \A_DOUT_TEMPR104[1] , 
        \A_DOUT_TEMPR104[0] }), .B_DOUT({nc11385, nc11386, nc11387, 
        nc11388, nc11389, nc11390, nc11391, nc11392, nc11393, nc11394, 
        nc11395, nc11396, nc11397, nc11398, nc11399, 
        \B_DOUT_TEMPR104[4] , \B_DOUT_TEMPR104[3] , 
        \B_DOUT_TEMPR104[2] , \B_DOUT_TEMPR104[1] , 
        \B_DOUT_TEMPR104[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[104][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1896 (.A(OR4_2972_Y), .B(OR4_837_Y), .C(OR4_484_Y), .D(
        OR4_1973_Y), .Y(OR4_1896_Y));
    OR4 OR4_817 (.A(OR4_373_Y), .B(OR4_2649_Y), .C(OR4_2381_Y), .D(
        OR4_1896_Y), .Y(OR4_817_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%48%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R48C6 (
        .A_DOUT({nc11400, nc11401, nc11402, nc11403, nc11404, nc11405, 
        nc11406, nc11407, nc11408, nc11409, nc11410, nc11411, nc11412, 
        nc11413, nc11414, \A_DOUT_TEMPR48[34] , \A_DOUT_TEMPR48[33] , 
        \A_DOUT_TEMPR48[32] , \A_DOUT_TEMPR48[31] , 
        \A_DOUT_TEMPR48[30] }), .B_DOUT({nc11415, nc11416, nc11417, 
        nc11418, nc11419, nc11420, nc11421, nc11422, nc11423, nc11424, 
        nc11425, nc11426, nc11427, nc11428, nc11429, 
        \B_DOUT_TEMPR48[34] , \B_DOUT_TEMPR48[33] , 
        \B_DOUT_TEMPR48[32] , \B_DOUT_TEMPR48[31] , 
        \B_DOUT_TEMPR48[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[48][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1419 (.A(\B_DOUT_TEMPR91[14] ), .B(\B_DOUT_TEMPR92[14] ), 
        .C(\B_DOUT_TEMPR93[14] ), .D(\B_DOUT_TEMPR94[14] ), .Y(
        OR4_1419_Y));
    OR4 OR4_1954 (.A(\A_DOUT_TEMPR83[28] ), .B(\A_DOUT_TEMPR84[28] ), 
        .C(\A_DOUT_TEMPR85[28] ), .D(\A_DOUT_TEMPR86[28] ), .Y(
        OR4_1954_Y));
    OR4 OR4_734 (.A(\B_DOUT_TEMPR107[10] ), .B(\B_DOUT_TEMPR108[10] ), 
        .C(\B_DOUT_TEMPR109[10] ), .D(\B_DOUT_TEMPR110[10] ), .Y(
        OR4_734_Y));
    OR4 OR4_2885 (.A(\B_DOUT_TEMPR75[11] ), .B(\B_DOUT_TEMPR76[11] ), 
        .C(\B_DOUT_TEMPR77[11] ), .D(\B_DOUT_TEMPR78[11] ), .Y(
        OR4_2885_Y));
    OR4 OR4_2945 (.A(\B_DOUT_TEMPR68[10] ), .B(\B_DOUT_TEMPR69[10] ), 
        .C(\B_DOUT_TEMPR70[10] ), .D(\B_DOUT_TEMPR71[10] ), .Y(
        OR4_2945_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%16%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R16C7 (
        .A_DOUT({nc11430, nc11431, nc11432, nc11433, nc11434, nc11435, 
        nc11436, nc11437, nc11438, nc11439, nc11440, nc11441, nc11442, 
        nc11443, nc11444, \A_DOUT_TEMPR16[39] , \A_DOUT_TEMPR16[38] , 
        \A_DOUT_TEMPR16[37] , \A_DOUT_TEMPR16[36] , 
        \A_DOUT_TEMPR16[35] }), .B_DOUT({nc11445, nc11446, nc11447, 
        nc11448, nc11449, nc11450, nc11451, nc11452, nc11453, nc11454, 
        nc11455, nc11456, nc11457, nc11458, nc11459, 
        \B_DOUT_TEMPR16[39] , \B_DOUT_TEMPR16[38] , 
        \B_DOUT_TEMPR16[37] , \B_DOUT_TEMPR16[36] , 
        \B_DOUT_TEMPR16[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%36%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R36C5 (
        .A_DOUT({nc11460, nc11461, nc11462, nc11463, nc11464, nc11465, 
        nc11466, nc11467, nc11468, nc11469, nc11470, nc11471, nc11472, 
        nc11473, nc11474, \A_DOUT_TEMPR36[29] , \A_DOUT_TEMPR36[28] , 
        \A_DOUT_TEMPR36[27] , \A_DOUT_TEMPR36[26] , 
        \A_DOUT_TEMPR36[25] }), .B_DOUT({nc11475, nc11476, nc11477, 
        nc11478, nc11479, nc11480, nc11481, nc11482, nc11483, nc11484, 
        nc11485, nc11486, nc11487, nc11488, nc11489, 
        \B_DOUT_TEMPR36[29] , \B_DOUT_TEMPR36[28] , 
        \B_DOUT_TEMPR36[27] , \B_DOUT_TEMPR36[26] , 
        \B_DOUT_TEMPR36[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1174 (.A(\B_DOUT_TEMPR99[2] ), .B(\B_DOUT_TEMPR100[2] ), 
        .C(\B_DOUT_TEMPR101[2] ), .D(\B_DOUT_TEMPR102[2] ), .Y(
        OR4_1174_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%39%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R39C5 (
        .A_DOUT({nc11490, nc11491, nc11492, nc11493, nc11494, nc11495, 
        nc11496, nc11497, nc11498, nc11499, nc11500, nc11501, nc11502, 
        nc11503, nc11504, \A_DOUT_TEMPR39[29] , \A_DOUT_TEMPR39[28] , 
        \A_DOUT_TEMPR39[27] , \A_DOUT_TEMPR39[26] , 
        \A_DOUT_TEMPR39[25] }), .B_DOUT({nc11505, nc11506, nc11507, 
        nc11508, nc11509, nc11510, nc11511, nc11512, nc11513, nc11514, 
        nc11515, nc11516, nc11517, nc11518, nc11519, 
        \B_DOUT_TEMPR39[29] , \B_DOUT_TEMPR39[28] , 
        \B_DOUT_TEMPR39[27] , \B_DOUT_TEMPR39[26] , 
        \B_DOUT_TEMPR39[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[39][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1956 (.A(OR4_1776_Y), .B(OR4_603_Y), .C(OR4_131_Y), .D(
        OR4_2206_Y), .Y(OR4_1956_Y));
    OR4 OR4_1642 (.A(\B_DOUT_TEMPR107[12] ), .B(\B_DOUT_TEMPR108[12] ), 
        .C(\B_DOUT_TEMPR109[12] ), .D(\B_DOUT_TEMPR110[12] ), .Y(
        OR4_1642_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_4 (.A(A_ADDR[16]), .B(A_ADDR[15]), .C(
        A_ADDR[14]), .Y(CFG3_4_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%69%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R69C3 (
        .A_DOUT({nc11520, nc11521, nc11522, nc11523, nc11524, nc11525, 
        nc11526, nc11527, nc11528, nc11529, nc11530, nc11531, nc11532, 
        nc11533, nc11534, \A_DOUT_TEMPR69[19] , \A_DOUT_TEMPR69[18] , 
        \A_DOUT_TEMPR69[17] , \A_DOUT_TEMPR69[16] , 
        \A_DOUT_TEMPR69[15] }), .B_DOUT({nc11535, nc11536, nc11537, 
        nc11538, nc11539, nc11540, nc11541, nc11542, nc11543, nc11544, 
        nc11545, nc11546, nc11547, nc11548, nc11549, 
        \B_DOUT_TEMPR69[19] , \B_DOUT_TEMPR69[18] , 
        \B_DOUT_TEMPR69[17] , \B_DOUT_TEMPR69[16] , 
        \B_DOUT_TEMPR69[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[69][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2649 (.A(OR4_1771_Y), .B(OR4_233_Y), .C(OR4_825_Y), .D(
        OR4_635_Y), .Y(OR4_2649_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%17%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R17C6 (
        .A_DOUT({nc11550, nc11551, nc11552, nc11553, nc11554, nc11555, 
        nc11556, nc11557, nc11558, nc11559, nc11560, nc11561, nc11562, 
        nc11563, nc11564, \A_DOUT_TEMPR17[34] , \A_DOUT_TEMPR17[33] , 
        \A_DOUT_TEMPR17[32] , \A_DOUT_TEMPR17[31] , 
        \A_DOUT_TEMPR17[30] }), .B_DOUT({nc11565, nc11566, nc11567, 
        nc11568, nc11569, nc11570, nc11571, nc11572, nc11573, nc11574, 
        nc11575, nc11576, nc11577, nc11578, nc11579, 
        \B_DOUT_TEMPR17[34] , \B_DOUT_TEMPR17[33] , 
        \B_DOUT_TEMPR17[32] , \B_DOUT_TEMPR17[31] , 
        \B_DOUT_TEMPR17[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_3007 (.A(\B_DOUT_TEMPR0[27] ), .B(\B_DOUT_TEMPR1[27] ), .C(
        \B_DOUT_TEMPR2[27] ), .D(\B_DOUT_TEMPR3[27] ), .Y(OR4_3007_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%81%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R81C4 (
        .A_DOUT({nc11580, nc11581, nc11582, nc11583, nc11584, nc11585, 
        nc11586, nc11587, nc11588, nc11589, nc11590, nc11591, nc11592, 
        nc11593, nc11594, \A_DOUT_TEMPR81[24] , \A_DOUT_TEMPR81[23] , 
        \A_DOUT_TEMPR81[22] , \A_DOUT_TEMPR81[21] , 
        \A_DOUT_TEMPR81[20] }), .B_DOUT({nc11595, nc11596, nc11597, 
        nc11598, nc11599, nc11600, nc11601, nc11602, nc11603, nc11604, 
        nc11605, nc11606, nc11607, nc11608, nc11609, 
        \B_DOUT_TEMPR81[24] , \B_DOUT_TEMPR81[23] , 
        \B_DOUT_TEMPR81[22] , \B_DOUT_TEMPR81[21] , 
        \B_DOUT_TEMPR81[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[81][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%99%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R99C7 (
        .A_DOUT({nc11610, nc11611, nc11612, nc11613, nc11614, nc11615, 
        nc11616, nc11617, nc11618, nc11619, nc11620, nc11621, nc11622, 
        nc11623, nc11624, \A_DOUT_TEMPR99[39] , \A_DOUT_TEMPR99[38] , 
        \A_DOUT_TEMPR99[37] , \A_DOUT_TEMPR99[36] , 
        \A_DOUT_TEMPR99[35] }), .B_DOUT({nc11625, nc11626, nc11627, 
        nc11628, nc11629, nc11630, nc11631, nc11632, nc11633, nc11634, 
        nc11635, nc11636, nc11637, nc11638, nc11639, 
        \B_DOUT_TEMPR99[39] , \B_DOUT_TEMPR99[38] , 
        \B_DOUT_TEMPR99[37] , \B_DOUT_TEMPR99[36] , 
        \B_DOUT_TEMPR99[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[99][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1942 (.A(\A_DOUT_TEMPR79[30] ), .B(\A_DOUT_TEMPR80[30] ), 
        .C(\A_DOUT_TEMPR81[30] ), .D(\A_DOUT_TEMPR82[30] ), .Y(
        OR4_1942_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%110%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R110C4 (
        .A_DOUT({nc11640, nc11641, nc11642, nc11643, nc11644, nc11645, 
        nc11646, nc11647, nc11648, nc11649, nc11650, nc11651, nc11652, 
        nc11653, nc11654, \A_DOUT_TEMPR110[24] , \A_DOUT_TEMPR110[23] , 
        \A_DOUT_TEMPR110[22] , \A_DOUT_TEMPR110[21] , 
        \A_DOUT_TEMPR110[20] }), .B_DOUT({nc11655, nc11656, nc11657, 
        nc11658, nc11659, nc11660, nc11661, nc11662, nc11663, nc11664, 
        nc11665, nc11666, nc11667, nc11668, nc11669, 
        \B_DOUT_TEMPR110[24] , \B_DOUT_TEMPR110[23] , 
        \B_DOUT_TEMPR110[22] , \B_DOUT_TEMPR110[21] , 
        \B_DOUT_TEMPR110[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[110][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_937 (.A(\A_DOUT_TEMPR91[0] ), .B(\A_DOUT_TEMPR92[0] ), .C(
        \A_DOUT_TEMPR93[0] ), .D(\A_DOUT_TEMPR94[0] ), .Y(OR4_937_Y));
    OR4 OR4_196 (.A(\B_DOUT_TEMPR4[30] ), .B(\B_DOUT_TEMPR5[30] ), .C(
        \B_DOUT_TEMPR6[30] ), .D(\B_DOUT_TEMPR7[30] ), .Y(OR4_196_Y));
    OR4 OR4_1260 (.A(\A_DOUT_TEMPR75[30] ), .B(\A_DOUT_TEMPR76[30] ), 
        .C(\A_DOUT_TEMPR77[30] ), .D(\A_DOUT_TEMPR78[30] ), .Y(
        OR4_1260_Y));
    OR4 OR4_1310 (.A(\B_DOUT_TEMPR68[16] ), .B(\B_DOUT_TEMPR69[16] ), 
        .C(\B_DOUT_TEMPR70[16] ), .D(\B_DOUT_TEMPR71[16] ), .Y(
        OR4_1310_Y));
    OR4 OR4_24 (.A(OR4_3020_Y), .B(OR4_1881_Y), .C(OR4_2512_Y), .D(
        OR4_1686_Y), .Y(OR4_24_Y));
    OR4 OR4_1417 (.A(\A_DOUT_TEMPR95[9] ), .B(\A_DOUT_TEMPR96[9] ), .C(
        \A_DOUT_TEMPR97[9] ), .D(\A_DOUT_TEMPR98[9] ), .Y(OR4_1417_Y));
    OR4 OR4_2527 (.A(OR4_1693_Y), .B(OR4_2654_Y), .C(OR4_1448_Y), .D(
        OR4_519_Y), .Y(OR4_2527_Y));
    OR4 OR4_2459 (.A(\A_DOUT_TEMPR64[1] ), .B(\A_DOUT_TEMPR65[1] ), .C(
        \A_DOUT_TEMPR66[1] ), .D(\A_DOUT_TEMPR67[1] ), .Y(OR4_2459_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%12%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R12C4 (
        .A_DOUT({nc11670, nc11671, nc11672, nc11673, nc11674, nc11675, 
        nc11676, nc11677, nc11678, nc11679, nc11680, nc11681, nc11682, 
        nc11683, nc11684, \A_DOUT_TEMPR12[24] , \A_DOUT_TEMPR12[23] , 
        \A_DOUT_TEMPR12[22] , \A_DOUT_TEMPR12[21] , 
        \A_DOUT_TEMPR12[20] }), .B_DOUT({nc11685, nc11686, nc11687, 
        nc11688, nc11689, nc11690, nc11691, nc11692, nc11693, nc11694, 
        nc11695, nc11696, nc11697, nc11698, nc11699, 
        \B_DOUT_TEMPR12[24] , \B_DOUT_TEMPR12[23] , 
        \B_DOUT_TEMPR12[22] , \B_DOUT_TEMPR12[21] , 
        \B_DOUT_TEMPR12[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_147 (.A(\B_DOUT_TEMPR28[1] ), .B(\B_DOUT_TEMPR29[1] ), .C(
        \B_DOUT_TEMPR30[1] ), .D(\B_DOUT_TEMPR31[1] ), .Y(OR4_147_Y));
    OR4 OR4_3020 (.A(OR4_1429_Y), .B(OR4_2222_Y), .C(OR2_31_Y), .D(
        \A_DOUT_TEMPR74[23] ), .Y(OR4_3020_Y));
    OR4 OR4_2660 (.A(\B_DOUT_TEMPR8[19] ), .B(\B_DOUT_TEMPR9[19] ), .C(
        \B_DOUT_TEMPR10[19] ), .D(\B_DOUT_TEMPR11[19] ), .Y(OR4_2660_Y)
        );
    OR4 OR4_604 (.A(\A_DOUT_TEMPR95[23] ), .B(\A_DOUT_TEMPR96[23] ), 
        .C(\A_DOUT_TEMPR97[23] ), .D(\A_DOUT_TEMPR98[23] ), .Y(
        OR4_604_Y));
    OR4 OR4_1790 (.A(\A_DOUT_TEMPR56[26] ), .B(\A_DOUT_TEMPR57[26] ), 
        .C(\A_DOUT_TEMPR58[26] ), .D(\A_DOUT_TEMPR59[26] ), .Y(
        OR4_1790_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%112%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R112C3 (
        .A_DOUT({nc11700, nc11701, nc11702, nc11703, nc11704, nc11705, 
        nc11706, nc11707, nc11708, nc11709, nc11710, nc11711, nc11712, 
        nc11713, nc11714, \A_DOUT_TEMPR112[19] , \A_DOUT_TEMPR112[18] , 
        \A_DOUT_TEMPR112[17] , \A_DOUT_TEMPR112[16] , 
        \A_DOUT_TEMPR112[15] }), .B_DOUT({nc11715, nc11716, nc11717, 
        nc11718, nc11719, nc11720, nc11721, nc11722, nc11723, nc11724, 
        nc11725, nc11726, nc11727, nc11728, nc11729, 
        \B_DOUT_TEMPR112[19] , \B_DOUT_TEMPR112[18] , 
        \B_DOUT_TEMPR112[17] , \B_DOUT_TEMPR112[16] , 
        \B_DOUT_TEMPR112[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[112][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2917 (.A(\A_DOUT_TEMPR44[26] ), .B(\A_DOUT_TEMPR45[26] ), 
        .C(\A_DOUT_TEMPR46[26] ), .D(\A_DOUT_TEMPR47[26] ), .Y(
        OR4_2917_Y));
    OR4 OR4_2068 (.A(\A_DOUT_TEMPR87[19] ), .B(\A_DOUT_TEMPR88[19] ), 
        .C(\A_DOUT_TEMPR89[19] ), .D(\A_DOUT_TEMPR90[19] ), .Y(
        OR4_2068_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%67%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R67C3 (
        .A_DOUT({nc11730, nc11731, nc11732, nc11733, nc11734, nc11735, 
        nc11736, nc11737, nc11738, nc11739, nc11740, nc11741, nc11742, 
        nc11743, nc11744, \A_DOUT_TEMPR67[19] , \A_DOUT_TEMPR67[18] , 
        \A_DOUT_TEMPR67[17] , \A_DOUT_TEMPR67[16] , 
        \A_DOUT_TEMPR67[15] }), .B_DOUT({nc11745, nc11746, nc11747, 
        nc11748, nc11749, nc11750, nc11751, nc11752, nc11753, nc11754, 
        nc11755, nc11756, nc11757, nc11758, nc11759, 
        \B_DOUT_TEMPR67[19] , \B_DOUT_TEMPR67[18] , 
        \B_DOUT_TEMPR67[17] , \B_DOUT_TEMPR67[16] , 
        \B_DOUT_TEMPR67[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[67][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1875 (.A(\A_DOUT_TEMPR56[36] ), .B(\A_DOUT_TEMPR57[36] ), 
        .C(\A_DOUT_TEMPR58[36] ), .D(\A_DOUT_TEMPR59[36] ), .Y(
        OR4_1875_Y));
    OR4 OR4_536 (.A(\B_DOUT_TEMPR95[19] ), .B(\B_DOUT_TEMPR96[19] ), 
        .C(\B_DOUT_TEMPR97[19] ), .D(\B_DOUT_TEMPR98[19] ), .Y(
        OR4_536_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%29%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R29C1 (
        .A_DOUT({nc11760, nc11761, nc11762, nc11763, nc11764, nc11765, 
        nc11766, nc11767, nc11768, nc11769, nc11770, nc11771, nc11772, 
        nc11773, nc11774, \A_DOUT_TEMPR29[9] , \A_DOUT_TEMPR29[8] , 
        \A_DOUT_TEMPR29[7] , \A_DOUT_TEMPR29[6] , \A_DOUT_TEMPR29[5] })
        , .B_DOUT({nc11775, nc11776, nc11777, nc11778, nc11779, 
        nc11780, nc11781, nc11782, nc11783, nc11784, nc11785, nc11786, 
        nc11787, nc11788, nc11789, \B_DOUT_TEMPR29[9] , 
        \B_DOUT_TEMPR29[8] , \B_DOUT_TEMPR29[7] , \B_DOUT_TEMPR29[6] , 
        \B_DOUT_TEMPR29[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%81%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R81C3 (
        .A_DOUT({nc11790, nc11791, nc11792, nc11793, nc11794, nc11795, 
        nc11796, nc11797, nc11798, nc11799, nc11800, nc11801, nc11802, 
        nc11803, nc11804, \A_DOUT_TEMPR81[19] , \A_DOUT_TEMPR81[18] , 
        \A_DOUT_TEMPR81[17] , \A_DOUT_TEMPR81[16] , 
        \A_DOUT_TEMPR81[15] }), .B_DOUT({nc11805, nc11806, nc11807, 
        nc11808, nc11809, nc11810, nc11811, nc11812, nc11813, nc11814, 
        nc11815, nc11816, nc11817, nc11818, nc11819, 
        \B_DOUT_TEMPR81[19] , \B_DOUT_TEMPR81[18] , 
        \B_DOUT_TEMPR81[17] , \B_DOUT_TEMPR81[16] , 
        \B_DOUT_TEMPR81[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[81][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%44%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R44C3 (
        .A_DOUT({nc11820, nc11821, nc11822, nc11823, nc11824, nc11825, 
        nc11826, nc11827, nc11828, nc11829, nc11830, nc11831, nc11832, 
        nc11833, nc11834, \A_DOUT_TEMPR44[19] , \A_DOUT_TEMPR44[18] , 
        \A_DOUT_TEMPR44[17] , \A_DOUT_TEMPR44[16] , 
        \A_DOUT_TEMPR44[15] }), .B_DOUT({nc11835, nc11836, nc11837, 
        nc11838, nc11839, nc11840, nc11841, nc11842, nc11843, nc11844, 
        nc11845, nc11846, nc11847, nc11848, nc11849, 
        \B_DOUT_TEMPR44[19] , \B_DOUT_TEMPR44[18] , 
        \B_DOUT_TEMPR44[17] , \B_DOUT_TEMPR44[16] , 
        \B_DOUT_TEMPR44[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[44][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1288 (.A(\B_DOUT_TEMPR20[36] ), .B(\B_DOUT_TEMPR21[36] ), 
        .C(\B_DOUT_TEMPR22[36] ), .D(\B_DOUT_TEMPR23[36] ), .Y(
        OR4_1288_Y));
    OR4 OR4_226 (.A(\A_DOUT_TEMPR16[6] ), .B(\A_DOUT_TEMPR17[6] ), .C(
        \A_DOUT_TEMPR18[6] ), .D(\A_DOUT_TEMPR19[6] ), .Y(OR4_226_Y));
    OR4 OR4_1366 (.A(\B_DOUT_TEMPR44[38] ), .B(\B_DOUT_TEMPR45[38] ), 
        .C(\B_DOUT_TEMPR46[38] ), .D(\B_DOUT_TEMPR47[38] ), .Y(
        OR4_1366_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%29%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R29C2 (
        .A_DOUT({nc11850, nc11851, nc11852, nc11853, nc11854, nc11855, 
        nc11856, nc11857, nc11858, nc11859, nc11860, nc11861, nc11862, 
        nc11863, nc11864, \A_DOUT_TEMPR29[14] , \A_DOUT_TEMPR29[13] , 
        \A_DOUT_TEMPR29[12] , \A_DOUT_TEMPR29[11] , 
        \A_DOUT_TEMPR29[10] }), .B_DOUT({nc11865, nc11866, nc11867, 
        nc11868, nc11869, nc11870, nc11871, nc11872, nc11873, nc11874, 
        nc11875, nc11876, nc11877, nc11878, nc11879, 
        \B_DOUT_TEMPR29[14] , \B_DOUT_TEMPR29[13] , 
        \B_DOUT_TEMPR29[12] , \B_DOUT_TEMPR29[11] , 
        \B_DOUT_TEMPR29[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2350 (.A(\B_DOUT_TEMPR28[31] ), .B(\B_DOUT_TEMPR29[31] ), 
        .C(\B_DOUT_TEMPR30[31] ), .D(\B_DOUT_TEMPR31[31] ), .Y(
        OR4_2350_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%25%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R25C1 (
        .A_DOUT({nc11880, nc11881, nc11882, nc11883, nc11884, nc11885, 
        nc11886, nc11887, nc11888, nc11889, nc11890, nc11891, nc11892, 
        nc11893, nc11894, \A_DOUT_TEMPR25[9] , \A_DOUT_TEMPR25[8] , 
        \A_DOUT_TEMPR25[7] , \A_DOUT_TEMPR25[6] , \A_DOUT_TEMPR25[5] })
        , .B_DOUT({nc11895, nc11896, nc11897, nc11898, nc11899, 
        nc11900, nc11901, nc11902, nc11903, nc11904, nc11905, nc11906, 
        nc11907, nc11908, nc11909, \B_DOUT_TEMPR25[9] , 
        \B_DOUT_TEMPR25[8] , \B_DOUT_TEMPR25[7] , \B_DOUT_TEMPR25[6] , 
        \B_DOUT_TEMPR25[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2457 (.A(\B_DOUT_TEMPR24[16] ), .B(\B_DOUT_TEMPR25[16] ), 
        .C(\B_DOUT_TEMPR26[16] ), .D(\B_DOUT_TEMPR27[16] ), .Y(
        OR4_2457_Y));
    OR4 OR4_593 (.A(OR4_1031_Y), .B(OR4_2574_Y), .C(OR4_352_Y), .D(
        OR4_2410_Y), .Y(OR4_593_Y));
    OR4 OR4_677 (.A(\A_DOUT_TEMPR103[4] ), .B(\A_DOUT_TEMPR104[4] ), 
        .C(\A_DOUT_TEMPR105[4] ), .D(\A_DOUT_TEMPR106[4] ), .Y(
        OR4_677_Y));
    OR4 OR4_2810 (.A(\B_DOUT_TEMPR107[21] ), .B(\B_DOUT_TEMPR108[21] ), 
        .C(\B_DOUT_TEMPR109[21] ), .D(\B_DOUT_TEMPR110[21] ), .Y(
        OR4_2810_Y));
    OR4 OR4_1397 (.A(OR4_1360_Y), .B(OR4_562_Y), .C(OR4_1271_Y), .D(
        OR4_1549_Y), .Y(OR4_1397_Y));
    OR4 OR4_1292 (.A(\B_DOUT_TEMPR56[37] ), .B(\B_DOUT_TEMPR57[37] ), 
        .C(\B_DOUT_TEMPR58[37] ), .D(\B_DOUT_TEMPR59[37] ), .Y(
        OR4_1292_Y));
    OR4 OR4_411 (.A(\B_DOUT_TEMPR107[39] ), .B(\B_DOUT_TEMPR108[39] ), 
        .C(\B_DOUT_TEMPR109[39] ), .D(\B_DOUT_TEMPR110[39] ), .Y(
        OR4_411_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%80%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R80C2 (
        .A_DOUT({nc11910, nc11911, nc11912, nc11913, nc11914, nc11915, 
        nc11916, nc11917, nc11918, nc11919, nc11920, nc11921, nc11922, 
        nc11923, nc11924, \A_DOUT_TEMPR80[14] , \A_DOUT_TEMPR80[13] , 
        \A_DOUT_TEMPR80[12] , \A_DOUT_TEMPR80[11] , 
        \A_DOUT_TEMPR80[10] }), .B_DOUT({nc11925, nc11926, nc11927, 
        nc11928, nc11929, nc11930, nc11931, nc11932, nc11933, nc11934, 
        nc11935, nc11936, nc11937, nc11938, nc11939, 
        \B_DOUT_TEMPR80[14] , \B_DOUT_TEMPR80[13] , 
        \B_DOUT_TEMPR80[12] , \B_DOUT_TEMPR80[11] , 
        \B_DOUT_TEMPR80[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[80][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2814 (.A(OR4_1167_Y), .B(OR4_155_Y), .C(OR4_375_Y), .D(
        OR4_170_Y), .Y(OR4_2814_Y));
    OR4 OR4_2164 (.A(OR4_587_Y), .B(OR4_1767_Y), .C(OR4_2844_Y), .D(
        OR4_2155_Y), .Y(OR4_2164_Y));
    OR4 OR4_1721 (.A(OR4_2088_Y), .B(OR4_3017_Y), .C(OR4_2662_Y), .D(
        OR4_1126_Y), .Y(OR4_1721_Y));
    OR4 OR4_1449 (.A(\B_DOUT_TEMPR79[36] ), .B(\B_DOUT_TEMPR80[36] ), 
        .C(\B_DOUT_TEMPR81[36] ), .D(\B_DOUT_TEMPR82[36] ), .Y(
        OR4_1449_Y));
    OR4 OR4_2698 (.A(\A_DOUT_TEMPR56[11] ), .B(\A_DOUT_TEMPR57[11] ), 
        .C(\A_DOUT_TEMPR58[11] ), .D(\A_DOUT_TEMPR59[11] ), .Y(
        OR4_2698_Y));
    OR4 OR4_2228 (.A(OR4_875_Y), .B(OR4_1839_Y), .C(OR4_2532_Y), .D(
        OR4_1174_Y), .Y(OR4_2228_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%70%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R70C0 (
        .A_DOUT({nc11940, nc11941, nc11942, nc11943, nc11944, nc11945, 
        nc11946, nc11947, nc11948, nc11949, nc11950, nc11951, nc11952, 
        nc11953, nc11954, \A_DOUT_TEMPR70[4] , \A_DOUT_TEMPR70[3] , 
        \A_DOUT_TEMPR70[2] , \A_DOUT_TEMPR70[1] , \A_DOUT_TEMPR70[0] })
        , .B_DOUT({nc11955, nc11956, nc11957, nc11958, nc11959, 
        nc11960, nc11961, nc11962, nc11963, nc11964, nc11965, nc11966, 
        nc11967, nc11968, nc11969, \B_DOUT_TEMPR70[4] , 
        \B_DOUT_TEMPR70[3] , \B_DOUT_TEMPR70[2] , \B_DOUT_TEMPR70[1] , 
        \B_DOUT_TEMPR70[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[70][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2047 (.A(\A_DOUT_TEMPR64[32] ), .B(\A_DOUT_TEMPR65[32] ), 
        .C(\A_DOUT_TEMPR66[32] ), .D(\A_DOUT_TEMPR67[32] ), .Y(
        OR4_2047_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%75%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R75C4 (
        .A_DOUT({nc11970, nc11971, nc11972, nc11973, nc11974, nc11975, 
        nc11976, nc11977, nc11978, nc11979, nc11980, nc11981, nc11982, 
        nc11983, nc11984, \A_DOUT_TEMPR75[24] , \A_DOUT_TEMPR75[23] , 
        \A_DOUT_TEMPR75[22] , \A_DOUT_TEMPR75[21] , 
        \A_DOUT_TEMPR75[20] }), .B_DOUT({nc11985, nc11986, nc11987, 
        nc11988, nc11989, nc11990, nc11991, nc11992, nc11993, nc11994, 
        nc11995, nc11996, nc11997, nc11998, nc11999, 
        \B_DOUT_TEMPR75[24] , \B_DOUT_TEMPR75[23] , 
        \B_DOUT_TEMPR75[22] , \B_DOUT_TEMPR75[21] , 
        \B_DOUT_TEMPR75[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[75][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2349 (.A(OR4_1750_Y), .B(OR4_2054_Y), .C(OR4_621_Y), .D(
        OR4_1534_Y), .Y(OR4_2349_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[27]  (.A(CFG3_20_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[27] ));
    OR4 OR4_2247 (.A(\A_DOUT_TEMPR68[33] ), .B(\A_DOUT_TEMPR69[33] ), 
        .C(\A_DOUT_TEMPR70[33] ), .D(\A_DOUT_TEMPR71[33] ), .Y(
        OR4_2247_Y));
    OR4 OR4_1494 (.A(\A_DOUT_TEMPR4[1] ), .B(\A_DOUT_TEMPR5[1] ), .C(
        \A_DOUT_TEMPR6[1] ), .D(\A_DOUT_TEMPR7[1] ), .Y(OR4_1494_Y));
    OR4 OR4_277 (.A(OR4_1384_Y), .B(OR4_2339_Y), .C(OR4_21_Y), .D(
        OR4_293_Y), .Y(OR4_277_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[29]  (.A(CFG3_6_Y), .B(CFG3_9_Y)
        , .Y(\BLKY2[29] ));
    OR4 OR4_867 (.A(OR4_1426_Y), .B(OR4_2777_Y), .C(OR4_2385_Y), .D(
        OR4_409_Y), .Y(OR4_867_Y));
    OR4 OR4_5 (.A(\A_DOUT_TEMPR111[3] ), .B(\A_DOUT_TEMPR112[3] ), .C(
        \A_DOUT_TEMPR113[3] ), .D(\A_DOUT_TEMPR114[3] ), .Y(OR4_5_Y));
    OR4 OR4_246 (.A(\A_DOUT_TEMPR115[1] ), .B(\A_DOUT_TEMPR116[1] ), 
        .C(\A_DOUT_TEMPR117[1] ), .D(\A_DOUT_TEMPR118[1] ), .Y(
        OR4_246_Y));
    OR4 OR4_607 (.A(OR4_2789_Y), .B(OR4_1296_Y), .C(OR4_2110_Y), .D(
        OR4_1157_Y), .Y(OR4_607_Y));
    OR4 OR4_1462 (.A(\A_DOUT_TEMPR40[28] ), .B(\A_DOUT_TEMPR41[28] ), 
        .C(\A_DOUT_TEMPR42[28] ), .D(\A_DOUT_TEMPR43[28] ), .Y(
        OR4_1462_Y));
    OR4 OR4_2940 (.A(OR4_1552_Y), .B(OR4_1865_Y), .C(OR4_1689_Y), .D(
        OR4_2196_Y), .Y(OR4_2940_Y));
    OR4 OR4_929 (.A(\B_DOUT_TEMPR75[13] ), .B(\B_DOUT_TEMPR76[13] ), 
        .C(\B_DOUT_TEMPR77[13] ), .D(\B_DOUT_TEMPR78[13] ), .Y(
        OR4_929_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[23]  (.A(CFG3_13_Y), .B(
        CFG3_3_Y), .Y(\BLKX2[23] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%27%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R27C5 (
        .A_DOUT({nc12000, nc12001, nc12002, nc12003, nc12004, nc12005, 
        nc12006, nc12007, nc12008, nc12009, nc12010, nc12011, nc12012, 
        nc12013, nc12014, \A_DOUT_TEMPR27[29] , \A_DOUT_TEMPR27[28] , 
        \A_DOUT_TEMPR27[27] , \A_DOUT_TEMPR27[26] , 
        \A_DOUT_TEMPR27[25] }), .B_DOUT({nc12015, nc12016, nc12017, 
        nc12018, nc12019, nc12020, nc12021, nc12022, nc12023, nc12024, 
        nc12025, nc12026, nc12027, nc12028, nc12029, 
        \B_DOUT_TEMPR27[29] , \B_DOUT_TEMPR27[28] , 
        \B_DOUT_TEMPR27[27] , \B_DOUT_TEMPR27[26] , 
        \B_DOUT_TEMPR27[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1340 (.A(\A_DOUT_TEMPR107[36] ), .B(\A_DOUT_TEMPR108[36] ), 
        .C(\A_DOUT_TEMPR109[36] ), .D(\A_DOUT_TEMPR110[36] ), .Y(
        OR4_1340_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[25]  (.A(CFG3_8_Y), .B(CFG3_9_Y)
        , .Y(\BLKY2[25] ));
    OR4 OR4_2688 (.A(\A_DOUT_TEMPR91[39] ), .B(\A_DOUT_TEMPR92[39] ), 
        .C(\A_DOUT_TEMPR93[39] ), .D(\A_DOUT_TEMPR94[39] ), .Y(
        OR4_2688_Y));
    OR4 OR4_1447 (.A(\B_DOUT_TEMPR56[24] ), .B(\B_DOUT_TEMPR57[24] ), 
        .C(\B_DOUT_TEMPR58[24] ), .D(\B_DOUT_TEMPR59[24] ), .Y(
        OR4_1447_Y));
    OR4 OR4_1468 (.A(OR4_1007_Y), .B(OR4_1298_Y), .C(OR4_942_Y), .D(
        OR4_1316_Y), .Y(OR4_1468_Y));
    OR4 OR4_2865 (.A(OR4_326_Y), .B(OR4_1168_Y), .C(OR4_199_Y), .D(
        OR4_145_Y), .Y(OR4_2865_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%66%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R66C5 (
        .A_DOUT({nc12030, nc12031, nc12032, nc12033, nc12034, nc12035, 
        nc12036, nc12037, nc12038, nc12039, nc12040, nc12041, nc12042, 
        nc12043, nc12044, \A_DOUT_TEMPR66[29] , \A_DOUT_TEMPR66[28] , 
        \A_DOUT_TEMPR66[27] , \A_DOUT_TEMPR66[26] , 
        \A_DOUT_TEMPR66[25] }), .B_DOUT({nc12045, nc12046, nc12047, 
        nc12048, nc12049, nc12050, nc12051, nc12052, nc12053, nc12054, 
        nc12055, nc12056, nc12057, nc12058, nc12059, 
        \B_DOUT_TEMPR66[29] , \B_DOUT_TEMPR66[28] , 
        \B_DOUT_TEMPR66[27] , \B_DOUT_TEMPR66[26] , 
        \B_DOUT_TEMPR66[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[66][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_654 (.A(\B_DOUT_TEMPR24[32] ), .B(\B_DOUT_TEMPR25[32] ), 
        .C(\B_DOUT_TEMPR26[32] ), .D(\B_DOUT_TEMPR27[32] ), .Y(
        OR4_654_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%69%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R69C5 (
        .A_DOUT({nc12060, nc12061, nc12062, nc12063, nc12064, nc12065, 
        nc12066, nc12067, nc12068, nc12069, nc12070, nc12071, nc12072, 
        nc12073, nc12074, \A_DOUT_TEMPR69[29] , \A_DOUT_TEMPR69[28] , 
        \A_DOUT_TEMPR69[27] , \A_DOUT_TEMPR69[26] , 
        \A_DOUT_TEMPR69[25] }), .B_DOUT({nc12075, nc12076, nc12077, 
        nc12078, nc12079, nc12080, nc12081, nc12082, nc12083, nc12084, 
        nc12085, nc12086, nc12087, nc12088, nc12089, 
        \B_DOUT_TEMPR69[29] , \B_DOUT_TEMPR69[28] , 
        \B_DOUT_TEMPR69[27] , \B_DOUT_TEMPR69[26] , 
        \B_DOUT_TEMPR69[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[69][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2039 (.A(OR4_569_Y), .B(OR4_2816_Y), .C(OR4_1760_Y), .D(
        OR4_2073_Y), .Y(OR4_2039_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[10]  (.A(CFG3_10_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[10] ));
    OR4 OR4_972 (.A(\A_DOUT_TEMPR28[17] ), .B(\A_DOUT_TEMPR29[17] ), 
        .C(\A_DOUT_TEMPR30[17] ), .D(\A_DOUT_TEMPR31[17] ), .Y(
        OR4_972_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%19%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R19C3 (
        .A_DOUT({nc12090, nc12091, nc12092, nc12093, nc12094, nc12095, 
        nc12096, nc12097, nc12098, nc12099, nc12100, nc12101, nc12102, 
        nc12103, nc12104, \A_DOUT_TEMPR19[19] , \A_DOUT_TEMPR19[18] , 
        \A_DOUT_TEMPR19[17] , \A_DOUT_TEMPR19[16] , 
        \A_DOUT_TEMPR19[15] }), .B_DOUT({nc12105, nc12106, nc12107, 
        nc12108, nc12109, nc12110, nc12111, nc12112, nc12113, nc12114, 
        nc12115, nc12116, nc12117, nc12118, nc12119, 
        \B_DOUT_TEMPR19[19] , \B_DOUT_TEMPR19[18] , 
        \B_DOUT_TEMPR19[17] , \B_DOUT_TEMPR19[16] , 
        \B_DOUT_TEMPR19[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_3019 (.A(\B_DOUT_TEMPR56[15] ), .B(\B_DOUT_TEMPR57[15] ), 
        .C(\B_DOUT_TEMPR58[15] ), .D(\B_DOUT_TEMPR59[15] ), .Y(
        OR4_3019_Y));
    OR4 OR4_1108 (.A(OR4_1046_Y), .B(OR4_1834_Y), .C(OR2_27_Y), .D(
        \A_DOUT_TEMPR74[22] ), .Y(OR4_1108_Y));
    OR4 OR4_175 (.A(OR4_433_Y), .B(OR4_1625_Y), .C(OR2_68_Y), .D(
        \A_DOUT_TEMPR74[10] ), .Y(OR4_175_Y));
    OR4 OR4_2539 (.A(\A_DOUT_TEMPR32[1] ), .B(\A_DOUT_TEMPR33[1] ), .C(
        \A_DOUT_TEMPR34[1] ), .D(\A_DOUT_TEMPR35[1] ), .Y(OR4_2539_Y));
    OR4 OR4_1039 (.A(\A_DOUT_TEMPR103[10] ), .B(\A_DOUT_TEMPR104[10] ), 
        .C(\A_DOUT_TEMPR105[10] ), .D(\A_DOUT_TEMPR106[10] ), .Y(
        OR4_1039_Y));
    OR4 OR4_1423 (.A(\A_DOUT_TEMPR56[24] ), .B(\A_DOUT_TEMPR57[24] ), 
        .C(\A_DOUT_TEMPR58[24] ), .D(\A_DOUT_TEMPR59[24] ), .Y(
        OR4_1423_Y));
    OR2 OR2_28 (.A(\A_DOUT_TEMPR72[37] ), .B(\A_DOUT_TEMPR73[37] ), .Y(
        OR2_28_Y));
    OR4 OR4_970 (.A(OR4_1907_Y), .B(OR4_1110_Y), .C(OR4_65_Y), .D(
        OR4_366_Y), .Y(OR4_970_Y));
    OR4 OR4_1539 (.A(\A_DOUT_TEMPR44[31] ), .B(\A_DOUT_TEMPR45[31] ), 
        .C(\A_DOUT_TEMPR46[31] ), .D(\A_DOUT_TEMPR47[31] ), .Y(
        OR4_1539_Y));
    OR4 OR4_2742 (.A(\A_DOUT_TEMPR36[35] ), .B(\A_DOUT_TEMPR37[35] ), 
        .C(\A_DOUT_TEMPR38[35] ), .D(\A_DOUT_TEMPR39[35] ), .Y(
        OR4_2742_Y));
    OR4 OR4_32 (.A(\A_DOUT_TEMPR24[29] ), .B(\A_DOUT_TEMPR25[29] ), .C(
        \A_DOUT_TEMPR26[29] ), .D(\A_DOUT_TEMPR27[29] ), .Y(OR4_32_Y));
    OR4 OR4_1560 (.A(\A_DOUT_TEMPR16[5] ), .B(\A_DOUT_TEMPR17[5] ), .C(
        \A_DOUT_TEMPR18[5] ), .D(\A_DOUT_TEMPR19[5] ), .Y(OR4_1560_Y));
    OR4 OR4_2332 (.A(\B_DOUT_TEMPR95[9] ), .B(\B_DOUT_TEMPR96[9] ), .C(
        \B_DOUT_TEMPR97[9] ), .D(\B_DOUT_TEMPR98[9] ), .Y(OR4_2332_Y));
    OR4 OR4_2102 (.A(OR4_1930_Y), .B(OR4_1868_Y), .C(OR4_2503_Y), .D(
        OR4_1678_Y), .Y(OR4_2102_Y));
    OR4 OR4_1803 (.A(\B_DOUT_TEMPR8[30] ), .B(\B_DOUT_TEMPR9[30] ), .C(
        \B_DOUT_TEMPR10[30] ), .D(\B_DOUT_TEMPR11[30] ), .Y(OR4_1803_Y)
        );
    OR4 OR4_1014 (.A(\B_DOUT_TEMPR48[39] ), .B(\B_DOUT_TEMPR49[39] ), 
        .C(\B_DOUT_TEMPR50[39] ), .D(\B_DOUT_TEMPR51[39] ), .Y(
        OR4_1014_Y));
    OR4 OR4_1016 (.A(\A_DOUT_TEMPR99[23] ), .B(\A_DOUT_TEMPR100[23] ), 
        .C(\A_DOUT_TEMPR101[23] ), .D(\A_DOUT_TEMPR102[23] ), .Y(
        OR4_1016_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%17%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R17C3 (
        .A_DOUT({nc12120, nc12121, nc12122, nc12123, nc12124, nc12125, 
        nc12126, nc12127, nc12128, nc12129, nc12130, nc12131, nc12132, 
        nc12133, nc12134, \A_DOUT_TEMPR17[19] , \A_DOUT_TEMPR17[18] , 
        \A_DOUT_TEMPR17[17] , \A_DOUT_TEMPR17[16] , 
        \A_DOUT_TEMPR17[15] }), .B_DOUT({nc12135, nc12136, nc12137, 
        nc12138, nc12139, nc12140, nc12141, nc12142, nc12143, nc12144, 
        nc12145, nc12146, nc12147, nc12148, nc12149, 
        \B_DOUT_TEMPR17[19] , \B_DOUT_TEMPR17[18] , 
        \B_DOUT_TEMPR17[17] , \B_DOUT_TEMPR17[16] , 
        \B_DOUT_TEMPR17[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%59%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R59C7 (
        .A_DOUT({nc12150, nc12151, nc12152, nc12153, nc12154, nc12155, 
        nc12156, nc12157, nc12158, nc12159, nc12160, nc12161, nc12162, 
        nc12163, nc12164, \A_DOUT_TEMPR59[39] , \A_DOUT_TEMPR59[38] , 
        \A_DOUT_TEMPR59[37] , \A_DOUT_TEMPR59[36] , 
        \A_DOUT_TEMPR59[35] }), .B_DOUT({nc12165, nc12166, nc12167, 
        nc12168, nc12169, nc12170, nc12171, nc12172, nc12173, nc12174, 
        nc12175, nc12176, nc12177, nc12178, nc12179, 
        \B_DOUT_TEMPR59[39] , \B_DOUT_TEMPR59[38] , 
        \B_DOUT_TEMPR59[37] , \B_DOUT_TEMPR59[36] , 
        \B_DOUT_TEMPR59[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[59][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_207 (.A(\A_DOUT_TEMPR111[17] ), .B(\A_DOUT_TEMPR112[17] ), 
        .C(\A_DOUT_TEMPR113[17] ), .D(\A_DOUT_TEMPR114[17] ), .Y(
        OR4_207_Y));
    OR4 OR4_1332 (.A(\A_DOUT_TEMPR103[2] ), .B(\A_DOUT_TEMPR104[2] ), 
        .C(\A_DOUT_TEMPR105[2] ), .D(\A_DOUT_TEMPR106[2] ), .Y(
        OR4_1332_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[26]  (.A(CFG3_10_Y), .B(
        CFG3_18_Y), .Y(\BLKX2[26] ));
    OR4 OR4_283 (.A(\B_DOUT_TEMPR48[12] ), .B(\B_DOUT_TEMPR49[12] ), 
        .C(\B_DOUT_TEMPR50[12] ), .D(\B_DOUT_TEMPR51[12] ), .Y(
        OR4_283_Y));
    OR4 OR4_1709 (.A(\A_DOUT_TEMPR64[21] ), .B(\A_DOUT_TEMPR65[21] ), 
        .C(\A_DOUT_TEMPR66[21] ), .D(\A_DOUT_TEMPR67[21] ), .Y(
        OR4_1709_Y));
    OR4 OR4_1678 (.A(\A_DOUT_TEMPR44[21] ), .B(\A_DOUT_TEMPR45[21] ), 
        .C(\A_DOUT_TEMPR46[21] ), .D(\A_DOUT_TEMPR47[21] ), .Y(
        OR4_1678_Y));
    OR2 OR2_5 (.A(\B_DOUT_TEMPR72[7] ), .B(\B_DOUT_TEMPR73[7] ), .Y(
        OR2_5_Y));
    OR4 OR4_381 (.A(\B_DOUT_TEMPR56[26] ), .B(\B_DOUT_TEMPR57[26] ), 
        .C(\B_DOUT_TEMPR58[26] ), .D(\B_DOUT_TEMPR59[26] ), .Y(
        OR4_381_Y));
    OR4 OR4_1294 (.A(\B_DOUT_TEMPR115[10] ), .B(\B_DOUT_TEMPR116[10] ), 
        .C(\B_DOUT_TEMPR117[10] ), .D(\B_DOUT_TEMPR118[10] ), .Y(
        OR4_1294_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%25%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R25C7 (
        .A_DOUT({nc12180, nc12181, nc12182, nc12183, nc12184, nc12185, 
        nc12186, nc12187, nc12188, nc12189, nc12190, nc12191, nc12192, 
        nc12193, nc12194, \A_DOUT_TEMPR25[39] , \A_DOUT_TEMPR25[38] , 
        \A_DOUT_TEMPR25[37] , \A_DOUT_TEMPR25[36] , 
        \A_DOUT_TEMPR25[35] }), .B_DOUT({nc12195, nc12196, nc12197, 
        nc12198, nc12199, nc12200, nc12201, nc12202, nc12203, nc12204, 
        nc12205, nc12206, nc12207, nc12208, nc12209, 
        \B_DOUT_TEMPR25[39] , \B_DOUT_TEMPR25[38] , 
        \B_DOUT_TEMPR25[37] , \B_DOUT_TEMPR25[36] , 
        \B_DOUT_TEMPR25[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[8]  (.A(CFG3_17_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[8] ));
    OR4 OR4_885 (.A(OR4_2760_Y), .B(OR4_82_Y), .C(OR4_833_Y), .D(
        OR4_1633_Y), .Y(OR4_885_Y));
    OR4 OR4_183 (.A(\A_DOUT_TEMPR87[35] ), .B(\A_DOUT_TEMPR88[35] ), 
        .C(\A_DOUT_TEMPR89[35] ), .D(\A_DOUT_TEMPR90[35] ), .Y(
        OR4_183_Y));
    OR4 OR4_2642 (.A(\A_DOUT_TEMPR83[13] ), .B(\A_DOUT_TEMPR84[13] ), 
        .C(\A_DOUT_TEMPR85[13] ), .D(\A_DOUT_TEMPR86[13] ), .Y(
        OR4_2642_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%84%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R84C6 (
        .A_DOUT({nc12210, nc12211, nc12212, nc12213, nc12214, nc12215, 
        nc12216, nc12217, nc12218, nc12219, nc12220, nc12221, nc12222, 
        nc12223, nc12224, \A_DOUT_TEMPR84[34] , \A_DOUT_TEMPR84[33] , 
        \A_DOUT_TEMPR84[32] , \A_DOUT_TEMPR84[31] , 
        \A_DOUT_TEMPR84[30] }), .B_DOUT({nc12225, nc12226, nc12227, 
        nc12228, nc12229, nc12230, nc12231, nc12232, nc12233, nc12234, 
        nc12235, nc12236, nc12237, nc12238, nc12239, 
        \B_DOUT_TEMPR84[34] , \B_DOUT_TEMPR84[33] , 
        \B_DOUT_TEMPR84[32] , \B_DOUT_TEMPR84[31] , 
        \B_DOUT_TEMPR84[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[84][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%78%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R78C6 (
        .A_DOUT({nc12240, nc12241, nc12242, nc12243, nc12244, nc12245, 
        nc12246, nc12247, nc12248, nc12249, nc12250, nc12251, nc12252, 
        nc12253, nc12254, \A_DOUT_TEMPR78[34] , \A_DOUT_TEMPR78[33] , 
        \A_DOUT_TEMPR78[32] , \A_DOUT_TEMPR78[31] , 
        \A_DOUT_TEMPR78[30] }), .B_DOUT({nc12255, nc12256, nc12257, 
        nc12258, nc12259, nc12260, nc12261, nc12262, nc12263, nc12264, 
        nc12265, nc12266, nc12267, nc12268, nc12269, 
        \B_DOUT_TEMPR78[34] , \B_DOUT_TEMPR78[33] , 
        \B_DOUT_TEMPR78[32] , \B_DOUT_TEMPR78[31] , 
        \B_DOUT_TEMPR78[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[78][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1313 (.A(\A_DOUT_TEMPR107[26] ), .B(\A_DOUT_TEMPR108[26] ), 
        .C(\A_DOUT_TEMPR109[26] ), .D(\A_DOUT_TEMPR110[26] ), .Y(
        OR4_1313_Y));
    OR4 OR4_902 (.A(OR4_267_Y), .B(OR4_1688_Y), .C(OR4_1210_Y), .D(
        OR4_294_Y), .Y(OR4_902_Y));
    OR4 OR4_1106 (.A(OR4_2459_Y), .B(OR4_863_Y), .C(OR2_9_Y), .D(
        \A_DOUT_TEMPR74[1] ), .Y(OR4_1106_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%42%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R42C6 (
        .A_DOUT({nc12270, nc12271, nc12272, nc12273, nc12274, nc12275, 
        nc12276, nc12277, nc12278, nc12279, nc12280, nc12281, nc12282, 
        nc12283, nc12284, \A_DOUT_TEMPR42[34] , \A_DOUT_TEMPR42[33] , 
        \A_DOUT_TEMPR42[32] , \A_DOUT_TEMPR42[31] , 
        \A_DOUT_TEMPR42[30] }), .B_DOUT({nc12285, nc12286, nc12287, 
        nc12288, nc12289, nc12290, nc12291, nc12292, nc12293, nc12294, 
        nc12295, nc12296, nc12297, nc12298, nc12299, 
        \B_DOUT_TEMPR42[34] , \B_DOUT_TEMPR42[33] , 
        \B_DOUT_TEMPR42[32] , \B_DOUT_TEMPR42[31] , 
        \B_DOUT_TEMPR42[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[42][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2942 (.A(OR4_1730_Y), .B(OR4_758_Y), .C(OR4_998_Y), .D(
        OR4_772_Y), .Y(OR4_2942_Y));
    OR4 OR4_105 (.A(OR4_1717_Y), .B(OR4_408_Y), .C(OR4_2306_Y), .D(
        OR4_2523_Y), .Y(OR4_105_Y));
    OR4 OR4_949 (.A(\B_DOUT_TEMPR24[29] ), .B(\B_DOUT_TEMPR25[29] ), 
        .C(\B_DOUT_TEMPR26[29] ), .D(\B_DOUT_TEMPR27[29] ), .Y(
        OR4_949_Y));
    OR4 OR4_1508 (.A(OR4_510_Y), .B(OR4_2755_Y), .C(OR4_1694_Y), .D(
        OR4_2009_Y), .Y(OR4_1508_Y));
    OR4 OR4_819 (.A(\A_DOUT_TEMPR32[4] ), .B(\A_DOUT_TEMPR33[4] ), .C(
        \A_DOUT_TEMPR34[4] ), .D(\A_DOUT_TEMPR35[4] ), .Y(OR4_819_Y));
    OR4 OR4_130 (.A(\A_DOUT_TEMPR64[27] ), .B(\A_DOUT_TEMPR65[27] ), 
        .C(\A_DOUT_TEMPR66[27] ), .D(\A_DOUT_TEMPR67[27] ), .Y(
        OR4_130_Y));
    OR4 OR4_1093 (.A(\A_DOUT_TEMPR79[13] ), .B(\A_DOUT_TEMPR80[13] ), 
        .C(\A_DOUT_TEMPR81[13] ), .D(\A_DOUT_TEMPR82[13] ), .Y(
        OR4_1093_Y));
    OR4 OR4_2315 (.A(\A_DOUT_TEMPR44[8] ), .B(\A_DOUT_TEMPR45[8] ), .C(
        \A_DOUT_TEMPR46[8] ), .D(\A_DOUT_TEMPR47[8] ), .Y(OR4_2315_Y));
    OR4 OR4_2054 (.A(\A_DOUT_TEMPR4[33] ), .B(\A_DOUT_TEMPR5[33] ), .C(
        \A_DOUT_TEMPR6[33] ), .D(\A_DOUT_TEMPR7[33] ), .Y(OR4_2054_Y));
    OR4 OR4_2535 (.A(\B_DOUT_TEMPR64[36] ), .B(\B_DOUT_TEMPR65[36] ), 
        .C(\B_DOUT_TEMPR66[36] ), .D(\B_DOUT_TEMPR67[36] ), .Y(
        OR4_2535_Y));
    OR4 OR4_2056 (.A(OR4_2451_Y), .B(OR4_363_Y), .C(OR4_857_Y), .D(
        OR4_1594_Y), .Y(OR4_2056_Y));
    OR4 OR4_900 (.A(\B_DOUT_TEMPR60[6] ), .B(\B_DOUT_TEMPR61[6] ), .C(
        \B_DOUT_TEMPR62[6] ), .D(\B_DOUT_TEMPR63[6] ), .Y(OR4_900_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%49%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R49C0 (
        .A_DOUT({nc12300, nc12301, nc12302, nc12303, nc12304, nc12305, 
        nc12306, nc12307, nc12308, nc12309, nc12310, nc12311, nc12312, 
        nc12313, nc12314, \A_DOUT_TEMPR49[4] , \A_DOUT_TEMPR49[3] , 
        \A_DOUT_TEMPR49[2] , \A_DOUT_TEMPR49[1] , \A_DOUT_TEMPR49[0] })
        , .B_DOUT({nc12315, nc12316, nc12317, nc12318, nc12319, 
        nc12320, nc12321, nc12322, nc12323, nc12324, nc12325, nc12326, 
        nc12327, nc12328, nc12329, \B_DOUT_TEMPR49[4] , 
        \B_DOUT_TEMPR49[3] , \B_DOUT_TEMPR49[2] , \B_DOUT_TEMPR49[1] , 
        \B_DOUT_TEMPR49[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2899 (.A(OR4_516_Y), .B(OR4_686_Y), .C(OR4_1386_Y), .D(
        OR4_1663_Y), .Y(OR4_2899_Y));
    OR4 OR4_1691 (.A(\B_DOUT_TEMPR32[39] ), .B(\B_DOUT_TEMPR33[39] ), 
        .C(\B_DOUT_TEMPR34[39] ), .D(\B_DOUT_TEMPR35[39] ), .Y(
        OR4_1691_Y));
    OR4 \OR4_A_DOUT[7]  (.A(OR4_945_Y), .B(OR4_974_Y), .C(OR4_1214_Y), 
        .D(OR4_2807_Y), .Y(A_DOUT[7]));
    OR4 OR4_1965 (.A(\B_DOUT_TEMPR12[32] ), .B(\B_DOUT_TEMPR13[32] ), 
        .C(\B_DOUT_TEMPR14[32] ), .D(\B_DOUT_TEMPR15[32] ), .Y(
        OR4_1965_Y));
    OR4 OR4_211 (.A(\A_DOUT_TEMPR107[37] ), .B(\A_DOUT_TEMPR108[37] ), 
        .C(\A_DOUT_TEMPR109[37] ), .D(\A_DOUT_TEMPR110[37] ), .Y(
        OR4_211_Y));
    OR4 OR4_811 (.A(OR4_646_Y), .B(OR4_2501_Y), .C(OR4_2040_Y), .D(
        OR4_1107_Y), .Y(OR4_811_Y));
    OR4 OR4_461 (.A(\B_DOUT_TEMPR83[7] ), .B(\B_DOUT_TEMPR84[7] ), .C(
        \B_DOUT_TEMPR85[7] ), .D(\B_DOUT_TEMPR86[7] ), .Y(OR4_461_Y));
    OR4 OR4_1535 (.A(OR4_160_Y), .B(OR4_490_Y), .C(OR4_306_Y), .D(
        OR4_851_Y), .Y(OR4_1535_Y));
    OR4 OR4_1793 (.A(\B_DOUT_TEMPR40[7] ), .B(\B_DOUT_TEMPR41[7] ), .C(
        \B_DOUT_TEMPR42[7] ), .D(\B_DOUT_TEMPR43[7] ), .Y(OR4_1793_Y));
    OR4 OR4_782 (.A(\B_DOUT_TEMPR60[28] ), .B(\B_DOUT_TEMPR61[28] ), 
        .C(\B_DOUT_TEMPR62[28] ), .D(\B_DOUT_TEMPR63[28] ), .Y(
        OR4_782_Y));
    OR4 OR4_61 (.A(\A_DOUT_TEMPR52[1] ), .B(\A_DOUT_TEMPR53[1] ), .C(
        \A_DOUT_TEMPR54[1] ), .D(\A_DOUT_TEMPR55[1] ), .Y(OR4_61_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%45%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R45C6 (
        .A_DOUT({nc12330, nc12331, nc12332, nc12333, nc12334, nc12335, 
        nc12336, nc12337, nc12338, nc12339, nc12340, nc12341, nc12342, 
        nc12343, nc12344, \A_DOUT_TEMPR45[34] , \A_DOUT_TEMPR45[33] , 
        \A_DOUT_TEMPR45[32] , \A_DOUT_TEMPR45[31] , 
        \A_DOUT_TEMPR45[30] }), .B_DOUT({nc12345, nc12346, nc12347, 
        nc12348, nc12349, nc12350, nc12351, nc12352, nc12353, nc12354, 
        nc12355, nc12356, nc12357, nc12358, nc12359, 
        \B_DOUT_TEMPR45[34] , \B_DOUT_TEMPR45[33] , 
        \B_DOUT_TEMPR45[32] , \B_DOUT_TEMPR45[31] , 
        \B_DOUT_TEMPR45[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_657 (.A(\A_DOUT_TEMPR40[29] ), .B(\A_DOUT_TEMPR41[29] ), 
        .C(\A_DOUT_TEMPR42[29] ), .D(\A_DOUT_TEMPR43[29] ), .Y(
        OR4_657_Y));
    OR4 \OR4_A_DOUT[35]  (.A(OR4_982_Y), .B(OR4_838_Y), .C(OR4_18_Y), 
        .D(OR4_624_Y), .Y(A_DOUT[35]));
    OR4 OR4_1582 (.A(\B_DOUT_TEMPR60[27] ), .B(\B_DOUT_TEMPR61[27] ), 
        .C(\B_DOUT_TEMPR62[27] ), .D(\B_DOUT_TEMPR63[27] ), .Y(
        OR4_1582_Y));
    OR4 OR4_638 (.A(\A_DOUT_TEMPR87[2] ), .B(\A_DOUT_TEMPR88[2] ), .C(
        \A_DOUT_TEMPR89[2] ), .D(\A_DOUT_TEMPR90[2] ), .Y(OR4_638_Y));
    OR4 OR4_1195 (.A(\A_DOUT_TEMPR8[23] ), .B(\A_DOUT_TEMPR9[23] ), .C(
        \A_DOUT_TEMPR10[23] ), .D(\A_DOUT_TEMPR11[23] ), .Y(OR4_1195_Y)
        );
    OR4 OR4_1669 (.A(\A_DOUT_TEMPR24[0] ), .B(\A_DOUT_TEMPR25[0] ), .C(
        \A_DOUT_TEMPR26[0] ), .D(\A_DOUT_TEMPR27[0] ), .Y(OR4_1669_Y));
    OR4 OR4_386 (.A(\A_DOUT_TEMPR20[26] ), .B(\A_DOUT_TEMPR21[26] ), 
        .C(\A_DOUT_TEMPR22[26] ), .D(\A_DOUT_TEMPR23[26] ), .Y(
        OR4_386_Y));
    OR4 OR4_34 (.A(\B_DOUT_TEMPR99[39] ), .B(\B_DOUT_TEMPR100[39] ), 
        .C(\B_DOUT_TEMPR101[39] ), .D(\B_DOUT_TEMPR102[39] ), .Y(
        OR4_34_Y));
    OR4 OR4_2191 (.A(\B_DOUT_TEMPR36[8] ), .B(\B_DOUT_TEMPR37[8] ), .C(
        \B_DOUT_TEMPR38[8] ), .D(\B_DOUT_TEMPR39[8] ), .Y(OR4_2191_Y));
    OR4 OR4_2353 (.A(\B_DOUT_TEMPR8[20] ), .B(\B_DOUT_TEMPR9[20] ), .C(
        \B_DOUT_TEMPR10[20] ), .D(\B_DOUT_TEMPR11[20] ), .Y(OR4_2353_Y)
        );
    OR4 OR4_82 (.A(\B_DOUT_TEMPR20[26] ), .B(\B_DOUT_TEMPR21[26] ), .C(
        \B_DOUT_TEMPR22[26] ), .D(\B_DOUT_TEMPR23[26] ), .Y(OR4_82_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%39%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R39C7 (
        .A_DOUT({nc12360, nc12361, nc12362, nc12363, nc12364, nc12365, 
        nc12366, nc12367, nc12368, nc12369, nc12370, nc12371, nc12372, 
        nc12373, nc12374, \A_DOUT_TEMPR39[39] , \A_DOUT_TEMPR39[38] , 
        \A_DOUT_TEMPR39[37] , \A_DOUT_TEMPR39[36] , 
        \A_DOUT_TEMPR39[35] }), .B_DOUT({nc12375, nc12376, nc12377, 
        nc12378, nc12379, nc12380, nc12381, nc12382, nc12383, nc12384, 
        nc12385, nc12386, nc12387, nc12388, nc12389, 
        \B_DOUT_TEMPR39[39] , \B_DOUT_TEMPR39[38] , 
        \B_DOUT_TEMPR39[37] , \B_DOUT_TEMPR39[36] , 
        \B_DOUT_TEMPR39[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[39][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2095 (.A(\A_DOUT_TEMPR107[4] ), .B(\A_DOUT_TEMPR108[4] ), 
        .C(\A_DOUT_TEMPR109[4] ), .D(\A_DOUT_TEMPR110[4] ), .Y(
        OR4_2095_Y));
    OR4 OR4_2889 (.A(\B_DOUT_TEMPR83[11] ), .B(\B_DOUT_TEMPR84[11] ), 
        .C(\B_DOUT_TEMPR85[11] ), .D(\B_DOUT_TEMPR86[11] ), .Y(
        OR4_2889_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%74%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R74C3 (
        .A_DOUT({nc12390, nc12391, nc12392, nc12393, nc12394, nc12395, 
        nc12396, nc12397, nc12398, nc12399, nc12400, nc12401, nc12402, 
        nc12403, nc12404, \A_DOUT_TEMPR74[19] , \A_DOUT_TEMPR74[18] , 
        \A_DOUT_TEMPR74[17] , \A_DOUT_TEMPR74[16] , 
        \A_DOUT_TEMPR74[15] }), .B_DOUT({nc12405, nc12406, nc12407, 
        nc12408, nc12409, nc12410, nc12411, nc12412, nc12413, nc12414, 
        nc12415, nc12416, nc12417, nc12418, nc12419, 
        \B_DOUT_TEMPR74[19] , \B_DOUT_TEMPR74[18] , 
        \B_DOUT_TEMPR74[17] , \B_DOUT_TEMPR74[16] , 
        \B_DOUT_TEMPR74[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[74][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_587 (.A(\A_DOUT_TEMPR103[18] ), .B(\A_DOUT_TEMPR104[18] ), 
        .C(\A_DOUT_TEMPR105[18] ), .D(\A_DOUT_TEMPR106[18] ), .Y(
        OR4_587_Y));
    OR4 OR4_694 (.A(\A_DOUT_TEMPR83[24] ), .B(\A_DOUT_TEMPR84[24] ), 
        .C(\A_DOUT_TEMPR85[24] ), .D(\A_DOUT_TEMPR86[24] ), .Y(
        OR4_694_Y));
    OR4 OR4_931 (.A(\A_DOUT_TEMPR28[32] ), .B(\A_DOUT_TEMPR29[32] ), 
        .C(\A_DOUT_TEMPR30[32] ), .D(\A_DOUT_TEMPR31[32] ), .Y(
        OR4_931_Y));
    OR4 OR4_1091 (.A(\A_DOUT_TEMPR99[25] ), .B(\A_DOUT_TEMPR100[25] ), 
        .C(\A_DOUT_TEMPR101[25] ), .D(\A_DOUT_TEMPR102[25] ), .Y(
        OR4_1091_Y));
    OR4 OR4_2938 (.A(\B_DOUT_TEMPR115[23] ), .B(\B_DOUT_TEMPR116[23] ), 
        .C(\B_DOUT_TEMPR117[23] ), .D(\B_DOUT_TEMPR118[23] ), .Y(
        OR4_2938_Y));
    OR4 OR4_1226 (.A(OR4_940_Y), .B(OR4_1297_Y), .C(OR4_1975_Y), .D(
        OR4_2256_Y), .Y(OR4_1226_Y));
    OR4 OR4_1938 (.A(\B_DOUT_TEMPR103[26] ), .B(\B_DOUT_TEMPR104[26] ), 
        .C(\B_DOUT_TEMPR105[26] ), .D(\B_DOUT_TEMPR106[26] ), .Y(
        OR4_1938_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%16%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R16C5 (
        .A_DOUT({nc12420, nc12421, nc12422, nc12423, nc12424, nc12425, 
        nc12426, nc12427, nc12428, nc12429, nc12430, nc12431, nc12432, 
        nc12433, nc12434, \A_DOUT_TEMPR16[29] , \A_DOUT_TEMPR16[28] , 
        \A_DOUT_TEMPR16[27] , \A_DOUT_TEMPR16[26] , 
        \A_DOUT_TEMPR16[25] }), .B_DOUT({nc12435, nc12436, nc12437, 
        nc12438, nc12439, nc12440, nc12441, nc12442, nc12443, nc12444, 
        nc12445, nc12446, nc12447, nc12448, nc12449, 
        \B_DOUT_TEMPR16[29] , \B_DOUT_TEMPR16[28] , 
        \B_DOUT_TEMPR16[27] , \B_DOUT_TEMPR16[26] , 
        \B_DOUT_TEMPR16[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%19%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R19C5 (
        .A_DOUT({nc12450, nc12451, nc12452, nc12453, nc12454, nc12455, 
        nc12456, nc12457, nc12458, nc12459, nc12460, nc12461, nc12462, 
        nc12463, nc12464, \A_DOUT_TEMPR19[29] , \A_DOUT_TEMPR19[28] , 
        \A_DOUT_TEMPR19[27] , \A_DOUT_TEMPR19[26] , 
        \A_DOUT_TEMPR19[25] }), .B_DOUT({nc12465, nc12466, nc12467, 
        nc12468, nc12469, nc12470, nc12471, nc12472, nc12473, nc12474, 
        nc12475, nc12476, nc12477, nc12478, nc12479, 
        \B_DOUT_TEMPR19[29] , \B_DOUT_TEMPR19[28] , 
        \B_DOUT_TEMPR19[27] , \B_DOUT_TEMPR19[26] , 
        \B_DOUT_TEMPR19[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2181 (.A(\B_DOUT_TEMPR12[0] ), .B(\B_DOUT_TEMPR13[0] ), .C(
        \B_DOUT_TEMPR14[0] ), .D(\B_DOUT_TEMPR15[0] ), .Y(OR4_2181_Y));
    OR4 OR4_2668 (.A(\B_DOUT_TEMPR103[15] ), .B(\B_DOUT_TEMPR104[15] ), 
        .C(\B_DOUT_TEMPR105[15] ), .D(\B_DOUT_TEMPR106[15] ), .Y(
        OR4_2668_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%27%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R27C2 (
        .A_DOUT({nc12480, nc12481, nc12482, nc12483, nc12484, nc12485, 
        nc12486, nc12487, nc12488, nc12489, nc12490, nc12491, nc12492, 
        nc12493, nc12494, \A_DOUT_TEMPR27[14] , \A_DOUT_TEMPR27[13] , 
        \A_DOUT_TEMPR27[12] , \A_DOUT_TEMPR27[11] , 
        \A_DOUT_TEMPR27[10] }), .B_DOUT({nc12495, nc12496, nc12497, 
        nc12498, nc12499, nc12500, nc12501, nc12502, nc12503, nc12504, 
        nc12505, nc12506, nc12507, nc12508, nc12509, 
        \B_DOUT_TEMPR27[14] , \B_DOUT_TEMPR27[13] , 
        \B_DOUT_TEMPR27[12] , \B_DOUT_TEMPR27[11] , 
        \B_DOUT_TEMPR27[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2897 (.A(OR4_54_Y), .B(OR4_1121_Y), .C(OR4_2833_Y), .D(
        OR4_1212_Y), .Y(OR4_2897_Y));
    OR4 OR4_1044 (.A(OR4_1714_Y), .B(OR4_1077_Y), .C(OR2_78_Y), .D(
        \B_DOUT_TEMPR74[3] ), .Y(OR4_1044_Y));
    OR4 OR4_1046 (.A(\A_DOUT_TEMPR64[22] ), .B(\A_DOUT_TEMPR65[22] ), 
        .C(\A_DOUT_TEMPR66[22] ), .D(\A_DOUT_TEMPR67[22] ), .Y(
        OR4_1046_Y));
    OR4 OR4_257 (.A(\A_DOUT_TEMPR52[22] ), .B(\A_DOUT_TEMPR53[22] ), 
        .C(\A_DOUT_TEMPR54[22] ), .D(\A_DOUT_TEMPR55[22] ), .Y(
        OR4_257_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%96%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R96C1 (
        .A_DOUT({nc12510, nc12511, nc12512, nc12513, nc12514, nc12515, 
        nc12516, nc12517, nc12518, nc12519, nc12520, nc12521, nc12522, 
        nc12523, nc12524, \A_DOUT_TEMPR96[9] , \A_DOUT_TEMPR96[8] , 
        \A_DOUT_TEMPR96[7] , \A_DOUT_TEMPR96[6] , \A_DOUT_TEMPR96[5] })
        , .B_DOUT({nc12525, nc12526, nc12527, nc12528, nc12529, 
        nc12530, nc12531, nc12532, nc12533, nc12534, nc12535, nc12536, 
        nc12537, nc12538, nc12539, \B_DOUT_TEMPR96[9] , 
        \B_DOUT_TEMPR96[8] , \B_DOUT_TEMPR96[7] , \B_DOUT_TEMPR96[6] , 
        \B_DOUT_TEMPR96[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[96][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2209 (.A(\A_DOUT_TEMPR83[30] ), .B(\A_DOUT_TEMPR84[30] ), 
        .C(\A_DOUT_TEMPR85[30] ), .D(\A_DOUT_TEMPR86[30] ), .Y(
        OR4_2209_Y));
    OR4 OR4_2085 (.A(OR4_181_Y), .B(OR4_2235_Y), .C(OR4_2455_Y), .D(
        OR4_2245_Y), .Y(OR4_2085_Y));
    OR4 OR4_317 (.A(OR4_864_Y), .B(OR4_765_Y), .C(OR4_2227_Y), .D(
        OR4_767_Y), .Y(OR4_317_Y));
    OR4 OR4_2522 (.A(\A_DOUT_TEMPR0[5] ), .B(\A_DOUT_TEMPR1[5] ), .C(
        \A_DOUT_TEMPR2[5] ), .D(\A_DOUT_TEMPR3[5] ), .Y(OR4_2522_Y));
    OR4 OR4_2449 (.A(\A_DOUT_TEMPR103[21] ), .B(\A_DOUT_TEMPR104[21] ), 
        .C(\A_DOUT_TEMPR105[21] ), .D(\A_DOUT_TEMPR106[21] ), .Y(
        OR4_2449_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_18 (.A(VCC), .B(A_ADDR[18]), .C(
        A_ADDR[17]), .Y(CFG3_18_Y));
    OR4 OR4_818 (.A(\B_DOUT_TEMPR24[17] ), .B(\B_DOUT_TEMPR25[17] ), 
        .C(\B_DOUT_TEMPR26[17] ), .D(\B_DOUT_TEMPR27[17] ), .Y(
        OR4_818_Y));
    OR4 OR4_611 (.A(\B_DOUT_TEMPR28[28] ), .B(\B_DOUT_TEMPR29[28] ), 
        .C(\B_DOUT_TEMPR30[28] ), .D(\B_DOUT_TEMPR31[28] ), .Y(
        OR4_611_Y));
    OR4 OR4_1504 (.A(\A_DOUT_TEMPR111[34] ), .B(\A_DOUT_TEMPR112[34] ), 
        .C(\A_DOUT_TEMPR113[34] ), .D(\A_DOUT_TEMPR114[34] ), .Y(
        OR4_1504_Y));
    OR4 OR4_1879 (.A(\B_DOUT_TEMPR75[3] ), .B(\B_DOUT_TEMPR76[3] ), .C(
        \B_DOUT_TEMPR77[3] ), .D(\B_DOUT_TEMPR78[3] ), .Y(OR4_1879_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%96%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R96C2 (
        .A_DOUT({nc12540, nc12541, nc12542, nc12543, nc12544, nc12545, 
        nc12546, nc12547, nc12548, nc12549, nc12550, nc12551, nc12552, 
        nc12553, nc12554, \A_DOUT_TEMPR96[14] , \A_DOUT_TEMPR96[13] , 
        \A_DOUT_TEMPR96[12] , \A_DOUT_TEMPR96[11] , 
        \A_DOUT_TEMPR96[10] }), .B_DOUT({nc12555, nc12556, nc12557, 
        nc12558, nc12559, nc12560, nc12561, nc12562, nc12563, nc12564, 
        nc12565, nc12566, nc12567, nc12568, nc12569, 
        \B_DOUT_TEMPR96[14] , \B_DOUT_TEMPR96[13] , 
        \B_DOUT_TEMPR96[12] , \B_DOUT_TEMPR96[11] , 
        \B_DOUT_TEMPR96[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[96][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1080 (.A(\B_DOUT_TEMPR79[3] ), .B(\B_DOUT_TEMPR80[3] ), .C(
        \B_DOUT_TEMPR81[3] ), .D(\B_DOUT_TEMPR82[3] ), .Y(OR4_1080_Y));
    OR4 OR4_952 (.A(\A_DOUT_TEMPR16[21] ), .B(\A_DOUT_TEMPR17[21] ), 
        .C(\A_DOUT_TEMPR18[21] ), .D(\A_DOUT_TEMPR19[21] ), .Y(
        OR4_952_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[18]  (.A(CFG3_10_Y), .B(
        CFG3_3_Y), .Y(\BLKX2[18] ));
    OR4 OR4_1343 (.A(OR4_2097_Y), .B(OR4_2089_Y), .C(OR4_1644_Y), .D(
        OR4_289_Y), .Y(OR4_1343_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%90%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R90C6 (
        .A_DOUT({nc12570, nc12571, nc12572, nc12573, nc12574, nc12575, 
        nc12576, nc12577, nc12578, nc12579, nc12580, nc12581, nc12582, 
        nc12583, nc12584, \A_DOUT_TEMPR90[34] , \A_DOUT_TEMPR90[33] , 
        \A_DOUT_TEMPR90[32] , \A_DOUT_TEMPR90[31] , 
        \A_DOUT_TEMPR90[30] }), .B_DOUT({nc12585, nc12586, nc12587, 
        nc12588, nc12589, nc12590, nc12591, nc12592, nc12593, nc12594, 
        nc12595, nc12596, nc12597, nc12598, nc12599, 
        \B_DOUT_TEMPR90[34] , \B_DOUT_TEMPR90[33] , 
        \B_DOUT_TEMPR90[32] , \B_DOUT_TEMPR90[31] , 
        \B_DOUT_TEMPR90[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[90][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_155 (.A(\A_DOUT_TEMPR91[11] ), .B(\A_DOUT_TEMPR92[11] ), 
        .C(\A_DOUT_TEMPR93[11] ), .D(\A_DOUT_TEMPR94[11] ), .Y(
        OR4_155_Y));
    OR4 OR4_2137 (.A(\B_DOUT_TEMPR24[4] ), .B(\B_DOUT_TEMPR25[4] ), .C(
        \B_DOUT_TEMPR26[4] ), .D(\B_DOUT_TEMPR27[4] ), .Y(OR4_2137_Y));
    OR4 OR4_934 (.A(\A_DOUT_TEMPR64[36] ), .B(\A_DOUT_TEMPR65[36] ), 
        .C(\A_DOUT_TEMPR66[36] ), .D(\A_DOUT_TEMPR67[36] ), .Y(
        OR4_934_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%90%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R90C5 (
        .A_DOUT({nc12600, nc12601, nc12602, nc12603, nc12604, nc12605, 
        nc12606, nc12607, nc12608, nc12609, nc12610, nc12611, nc12612, 
        nc12613, nc12614, \A_DOUT_TEMPR90[29] , \A_DOUT_TEMPR90[28] , 
        \A_DOUT_TEMPR90[27] , \A_DOUT_TEMPR90[26] , 
        \A_DOUT_TEMPR90[25] }), .B_DOUT({nc12615, nc12616, nc12617, 
        nc12618, nc12619, nc12620, nc12621, nc12622, nc12623, nc12624, 
        nc12625, nc12626, nc12627, nc12628, nc12629, 
        \B_DOUT_TEMPR90[29] , \B_DOUT_TEMPR90[28] , 
        \B_DOUT_TEMPR90[27] , \B_DOUT_TEMPR90[26] , 
        \B_DOUT_TEMPR90[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[90][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_41 (.A(\A_DOUT_TEMPR32[13] ), .B(\A_DOUT_TEMPR33[13] ), .C(
        \A_DOUT_TEMPR34[13] ), .D(\A_DOUT_TEMPR35[13] ), .Y(OR4_41_Y));
    OR4 OR4_2634 (.A(\B_DOUT_TEMPR91[12] ), .B(\B_DOUT_TEMPR92[12] ), 
        .C(\B_DOUT_TEMPR93[12] ), .D(\B_DOUT_TEMPR94[12] ), .Y(
        OR4_2634_Y));
    OR4 \OR4_A_DOUT[9]  (.A(OR4_2511_Y), .B(OR4_1162_Y), .C(OR4_1054_Y)
        , .D(OR4_2616_Y), .Y(A_DOUT[9]));
    OR4 OR4_2887 (.A(\A_DOUT_TEMPR0[1] ), .B(\A_DOUT_TEMPR1[1] ), .C(
        \A_DOUT_TEMPR2[1] ), .D(\A_DOUT_TEMPR3[1] ), .Y(OR4_2887_Y));
    OR4 OR4_84 (.A(\A_DOUT_TEMPR52[25] ), .B(\A_DOUT_TEMPR53[25] ), .C(
        \A_DOUT_TEMPR54[25] ), .D(\A_DOUT_TEMPR55[25] ), .Y(OR4_84_Y));
    OR4 OR4_950 (.A(\B_DOUT_TEMPR83[20] ), .B(\B_DOUT_TEMPR84[20] ), 
        .C(\B_DOUT_TEMPR85[20] ), .D(\B_DOUT_TEMPR86[20] ), .Y(
        OR4_950_Y));
    OR4 OR4_1826 (.A(\A_DOUT_TEMPR48[3] ), .B(\A_DOUT_TEMPR49[3] ), .C(
        \A_DOUT_TEMPR50[3] ), .D(\A_DOUT_TEMPR51[3] ), .Y(OR4_1826_Y));
    OR4 OR4_2340 (.A(\B_DOUT_TEMPR60[3] ), .B(\B_DOUT_TEMPR61[3] ), .C(
        \B_DOUT_TEMPR62[3] ), .D(\B_DOUT_TEMPR63[3] ), .Y(OR4_2340_Y));
    OR4 OR4_1137 (.A(OR4_2819_Y), .B(OR4_52_Y), .C(OR4_2565_Y), .D(
        OR4_616_Y), .Y(OR4_1137_Y));
    OR4 OR4_414 (.A(\A_DOUT_TEMPR44[14] ), .B(\A_DOUT_TEMPR45[14] ), 
        .C(\A_DOUT_TEMPR46[14] ), .D(\A_DOUT_TEMPR47[14] ), .Y(
        OR4_414_Y));
    OR4 OR4_1171 (.A(\B_DOUT_TEMPR20[10] ), .B(\B_DOUT_TEMPR21[10] ), 
        .C(\B_DOUT_TEMPR22[10] ), .D(\B_DOUT_TEMPR23[10] ), .Y(
        OR4_1171_Y));
    OR4 OR4_2447 (.A(\A_DOUT_TEMPR64[33] ), .B(\A_DOUT_TEMPR65[33] ), 
        .C(\A_DOUT_TEMPR66[33] ), .D(\A_DOUT_TEMPR67[33] ), .Y(
        OR4_2447_Y));
    OR4 OR4_1634 (.A(\B_DOUT_TEMPR103[13] ), .B(\B_DOUT_TEMPR104[13] ), 
        .C(\B_DOUT_TEMPR105[13] ), .D(\B_DOUT_TEMPR106[13] ), .Y(
        OR4_1634_Y));
    OR4 OR4_1067 (.A(\B_DOUT_TEMPR115[5] ), .B(\B_DOUT_TEMPR116[5] ), 
        .C(\B_DOUT_TEMPR117[5] ), .D(\B_DOUT_TEMPR118[5] ), .Y(
        OR4_1067_Y));
    OR4 OR4_1075 (.A(\B_DOUT_TEMPR40[38] ), .B(\B_DOUT_TEMPR41[38] ), 
        .C(\B_DOUT_TEMPR42[38] ), .D(\B_DOUT_TEMPR43[38] ), .Y(
        OR4_1075_Y));
    OR4 OR4_1369 (.A(\B_DOUT_TEMPR8[12] ), .B(\B_DOUT_TEMPR9[12] ), .C(
        \B_DOUT_TEMPR10[12] ), .D(\B_DOUT_TEMPR11[12] ), .Y(OR4_1369_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%104%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R104C6 (
        .A_DOUT({nc12630, nc12631, nc12632, nc12633, nc12634, nc12635, 
        nc12636, nc12637, nc12638, nc12639, nc12640, nc12641, nc12642, 
        nc12643, nc12644, \A_DOUT_TEMPR104[34] , \A_DOUT_TEMPR104[33] , 
        \A_DOUT_TEMPR104[32] , \A_DOUT_TEMPR104[31] , 
        \A_DOUT_TEMPR104[30] }), .B_DOUT({nc12645, nc12646, nc12647, 
        nc12648, nc12649, nc12650, nc12651, nc12652, nc12653, nc12654, 
        nc12655, nc12656, nc12657, nc12658, nc12659, 
        \B_DOUT_TEMPR104[34] , \B_DOUT_TEMPR104[33] , 
        \B_DOUT_TEMPR104[32] , \B_DOUT_TEMPR104[31] , 
        \B_DOUT_TEMPR104[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[104][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1267 (.A(\B_DOUT_TEMPR24[25] ), .B(\B_DOUT_TEMPR25[25] ), 
        .C(\B_DOUT_TEMPR26[25] ), .D(\B_DOUT_TEMPR27[25] ), .Y(
        OR4_1267_Y));
    OR4 \OR4_A_DOUT[11]  (.A(OR4_486_Y), .B(OR4_75_Y), .C(OR4_2814_Y), 
        .D(OR4_1718_Y), .Y(A_DOUT[11]));
    OR4 OR4_1201 (.A(OR4_1647_Y), .B(OR4_2472_Y), .C(OR4_1536_Y), .D(
        OR4_2992_Y), .Y(OR4_1201_Y));
    OR4 OR4_869 (.A(\B_DOUT_TEMPR64[31] ), .B(\B_DOUT_TEMPR65[31] ), 
        .C(\B_DOUT_TEMPR66[31] ), .D(\B_DOUT_TEMPR67[31] ), .Y(
        OR4_869_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%7%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R7C2 (
        .A_DOUT({nc12660, nc12661, nc12662, nc12663, nc12664, nc12665, 
        nc12666, nc12667, nc12668, nc12669, nc12670, nc12671, nc12672, 
        nc12673, nc12674, \A_DOUT_TEMPR7[14] , \A_DOUT_TEMPR7[13] , 
        \A_DOUT_TEMPR7[12] , \A_DOUT_TEMPR7[11] , \A_DOUT_TEMPR7[10] })
        , .B_DOUT({nc12675, nc12676, nc12677, nc12678, nc12679, 
        nc12680, nc12681, nc12682, nc12683, nc12684, nc12685, nc12686, 
        nc12687, nc12688, nc12689, \B_DOUT_TEMPR7[14] , 
        \B_DOUT_TEMPR7[13] , \B_DOUT_TEMPR7[12] , \B_DOUT_TEMPR7[11] , 
        \B_DOUT_TEMPR7[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_697 (.A(\B_DOUT_TEMPR115[18] ), .B(\B_DOUT_TEMPR116[18] ), 
        .C(\B_DOUT_TEMPR117[18] ), .D(\B_DOUT_TEMPR118[18] ), .Y(
        OR4_697_Y));
    OR4 OR4_786 (.A(\B_DOUT_TEMPR48[23] ), .B(\B_DOUT_TEMPR49[23] ), 
        .C(\B_DOUT_TEMPR50[23] ), .D(\B_DOUT_TEMPR51[23] ), .Y(
        OR4_786_Y));
    OR4 OR4_1960 (.A(\B_DOUT_TEMPR44[5] ), .B(\B_DOUT_TEMPR45[5] ), .C(
        \B_DOUT_TEMPR46[5] ), .D(\B_DOUT_TEMPR47[5] ), .Y(OR4_1960_Y));
    OR4 OR4_2020 (.A(\A_DOUT_TEMPR64[2] ), .B(\A_DOUT_TEMPR65[2] ), .C(
        \A_DOUT_TEMPR66[2] ), .D(\A_DOUT_TEMPR67[2] ), .Y(OR4_2020_Y));
    OR4 OR4_261 (.A(\B_DOUT_TEMPR79[2] ), .B(\B_DOUT_TEMPR80[2] ), .C(
        \B_DOUT_TEMPR81[2] ), .D(\B_DOUT_TEMPR82[2] ), .Y(OR4_261_Y));
    OR4 OR4_861 (.A(\B_DOUT_TEMPR107[33] ), .B(\B_DOUT_TEMPR108[33] ), 
        .C(\B_DOUT_TEMPR109[33] ), .D(\B_DOUT_TEMPR110[33] ), .Y(
        OR4_861_Y));
    OR4 OR4_1486 (.A(OR4_2656_Y), .B(OR4_2000_Y), .C(OR4_2643_Y), .D(
        OR4_1813_Y), .Y(OR4_1486_Y));
    OR4 OR4_1877 (.A(\A_DOUT_TEMPR60[33] ), .B(\A_DOUT_TEMPR61[33] ), 
        .C(\A_DOUT_TEMPR62[33] ), .D(\A_DOUT_TEMPR63[33] ), .Y(
        OR4_1877_Y));
    OR4 OR4_1720 (.A(\A_DOUT_TEMPR103[23] ), .B(\A_DOUT_TEMPR104[23] ), 
        .C(\A_DOUT_TEMPR105[23] ), .D(\A_DOUT_TEMPR106[23] ), .Y(
        OR4_1720_Y));
    OR4 OR4_66 (.A(\B_DOUT_TEMPR91[7] ), .B(\B_DOUT_TEMPR92[7] ), .C(
        \B_DOUT_TEMPR93[7] ), .D(\B_DOUT_TEMPR94[7] ), .Y(OR4_66_Y));
    OR4 OR4_3004 (.A(\B_DOUT_TEMPR103[31] ), .B(\B_DOUT_TEMPR104[31] ), 
        .C(\B_DOUT_TEMPR105[31] ), .D(\B_DOUT_TEMPR106[31] ), .Y(
        OR4_3004_Y));
    OR4 \OR4_A_DOUT[5]  (.A(OR4_1956_Y), .B(OR4_2665_Y), .C(OR4_2404_Y)
        , .D(OR4_1687_Y), .Y(A_DOUT[5]));
    OR4 OR4_3006 (.A(OR4_2936_Y), .B(OR4_655_Y), .C(OR4_216_Y), .D(
        OR4_1898_Y), .Y(OR4_3006_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%88%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R88C0 (
        .A_DOUT({nc12690, nc12691, nc12692, nc12693, nc12694, nc12695, 
        nc12696, nc12697, nc12698, nc12699, nc12700, nc12701, nc12702, 
        nc12703, nc12704, \A_DOUT_TEMPR88[4] , \A_DOUT_TEMPR88[3] , 
        \A_DOUT_TEMPR88[2] , \A_DOUT_TEMPR88[1] , \A_DOUT_TEMPR88[0] })
        , .B_DOUT({nc12705, nc12706, nc12707, nc12708, nc12709, 
        nc12710, nc12711, nc12712, nc12713, nc12714, nc12715, nc12716, 
        nc12717, nc12718, nc12719, \B_DOUT_TEMPR88[4] , 
        \B_DOUT_TEMPR88[3] , \B_DOUT_TEMPR88[2] , \B_DOUT_TEMPR88[1] , 
        \B_DOUT_TEMPR88[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[88][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%69%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R69C7 (
        .A_DOUT({nc12720, nc12721, nc12722, nc12723, nc12724, nc12725, 
        nc12726, nc12727, nc12728, nc12729, nc12730, nc12731, nc12732, 
        nc12733, nc12734, \A_DOUT_TEMPR69[39] , \A_DOUT_TEMPR69[38] , 
        \A_DOUT_TEMPR69[37] , \A_DOUT_TEMPR69[36] , 
        \A_DOUT_TEMPR69[35] }), .B_DOUT({nc12735, nc12736, nc12737, 
        nc12738, nc12739, nc12740, nc12741, nc12742, nc12743, nc12744, 
        nc12745, nc12746, nc12747, nc12748, nc12749, 
        \B_DOUT_TEMPR69[39] , \B_DOUT_TEMPR69[38] , 
        \B_DOUT_TEMPR69[37] , \B_DOUT_TEMPR69[36] , 
        \B_DOUT_TEMPR69[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[69][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%45%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R45C2 (
        .A_DOUT({nc12750, nc12751, nc12752, nc12753, nc12754, nc12755, 
        nc12756, nc12757, nc12758, nc12759, nc12760, nc12761, nc12762, 
        nc12763, nc12764, \A_DOUT_TEMPR45[14] , \A_DOUT_TEMPR45[13] , 
        \A_DOUT_TEMPR45[12] , \A_DOUT_TEMPR45[11] , 
        \A_DOUT_TEMPR45[10] }), .B_DOUT({nc12765, nc12766, nc12767, 
        nc12768, nc12769, nc12770, nc12771, nc12772, nc12773, nc12774, 
        nc12775, nc12776, nc12777, nc12778, nc12779, 
        \B_DOUT_TEMPR45[14] , \B_DOUT_TEMPR45[13] , 
        \B_DOUT_TEMPR45[12] , \B_DOUT_TEMPR45[11] , 
        \B_DOUT_TEMPR45[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1785 (.A(OR4_1036_Y), .B(OR4_1974_Y), .C(OR4_1276_Y), .D(
        OR4_988_Y), .Y(OR4_1785_Y));
    OR4 OR4_1762 (.A(\A_DOUT_TEMPR48[8] ), .B(\A_DOUT_TEMPR49[8] ), .C(
        \A_DOUT_TEMPR50[8] ), .D(\A_DOUT_TEMPR51[8] ), .Y(OR4_1762_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%1%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R1C6 (
        .A_DOUT({nc12780, nc12781, nc12782, nc12783, nc12784, nc12785, 
        nc12786, nc12787, nc12788, nc12789, nc12790, nc12791, nc12792, 
        nc12793, nc12794, \A_DOUT_TEMPR1[34] , \A_DOUT_TEMPR1[33] , 
        \A_DOUT_TEMPR1[32] , \A_DOUT_TEMPR1[31] , \A_DOUT_TEMPR1[30] })
        , .B_DOUT({nc12795, nc12796, nc12797, nc12798, nc12799, 
        nc12800, nc12801, nc12802, nc12803, nc12804, nc12805, nc12806, 
        nc12807, nc12808, nc12809, \B_DOUT_TEMPR1[34] , 
        \B_DOUT_TEMPR1[33] , \B_DOUT_TEMPR1[32] , \B_DOUT_TEMPR1[31] , 
        \B_DOUT_TEMPR1[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_581 (.A(\B_DOUT_TEMPR79[17] ), .B(\B_DOUT_TEMPR80[17] ), 
        .C(\B_DOUT_TEMPR81[17] ), .D(\B_DOUT_TEMPR82[17] ), .Y(
        OR4_581_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%116%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R116C2 (
        .A_DOUT({nc12810, nc12811, nc12812, nc12813, nc12814, nc12815, 
        nc12816, nc12817, nc12818, nc12819, nc12820, nc12821, nc12822, 
        nc12823, nc12824, \A_DOUT_TEMPR116[14] , \A_DOUT_TEMPR116[13] , 
        \A_DOUT_TEMPR116[12] , \A_DOUT_TEMPR116[11] , 
        \A_DOUT_TEMPR116[10] }), .B_DOUT({nc12825, nc12826, nc12827, 
        nc12828, nc12829, nc12830, nc12831, nc12832, nc12833, nc12834, 
        nc12835, nc12836, nc12837, nc12838, nc12839, 
        \B_DOUT_TEMPR116[14] , \B_DOUT_TEMPR116[13] , 
        \B_DOUT_TEMPR116[12] , \B_DOUT_TEMPR116[11] , 
        \B_DOUT_TEMPR116[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[116][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_588 (.A(\B_DOUT_TEMPR16[12] ), .B(\B_DOUT_TEMPR17[12] ), 
        .C(\B_DOUT_TEMPR18[12] ), .D(\B_DOUT_TEMPR19[12] ), .Y(
        OR4_588_Y));
    OR4 OR4_2869 (.A(\B_DOUT_TEMPR87[0] ), .B(\B_DOUT_TEMPR88[0] ), .C(
        \B_DOUT_TEMPR89[0] ), .D(\B_DOUT_TEMPR90[0] ), .Y(OR4_2869_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%109%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R109C1 (
        .A_DOUT({nc12840, nc12841, nc12842, nc12843, nc12844, nc12845, 
        nc12846, nc12847, nc12848, nc12849, nc12850, nc12851, nc12852, 
        nc12853, nc12854, \A_DOUT_TEMPR109[9] , \A_DOUT_TEMPR109[8] , 
        \A_DOUT_TEMPR109[7] , \A_DOUT_TEMPR109[6] , 
        \A_DOUT_TEMPR109[5] }), .B_DOUT({nc12855, nc12856, nc12857, 
        nc12858, nc12859, nc12860, nc12861, nc12862, nc12863, nc12864, 
        nc12865, nc12866, nc12867, nc12868, nc12869, 
        \B_DOUT_TEMPR109[9] , \B_DOUT_TEMPR109[8] , 
        \B_DOUT_TEMPR109[7] , \B_DOUT_TEMPR109[6] , 
        \B_DOUT_TEMPR109[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[109][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%98%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R98C5 (
        .A_DOUT({nc12870, nc12871, nc12872, nc12873, nc12874, nc12875, 
        nc12876, nc12877, nc12878, nc12879, nc12880, nc12881, nc12882, 
        nc12883, nc12884, \A_DOUT_TEMPR98[29] , \A_DOUT_TEMPR98[28] , 
        \A_DOUT_TEMPR98[27] , \A_DOUT_TEMPR98[26] , 
        \A_DOUT_TEMPR98[25] }), .B_DOUT({nc12885, nc12886, nc12887, 
        nc12888, nc12889, nc12890, nc12891, nc12892, nc12893, nc12894, 
        nc12895, nc12896, nc12897, nc12898, nc12899, 
        \B_DOUT_TEMPR98[29] , \B_DOUT_TEMPR98[28] , 
        \B_DOUT_TEMPR98[27] , \B_DOUT_TEMPR98[26] , 
        \B_DOUT_TEMPR98[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[98][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_73 (.A(\B_DOUT_TEMPR72[35] ), .B(\B_DOUT_TEMPR73[35] ), .Y(
        OR2_73_Y));
    OR4 OR4_297 (.A(OR4_909_Y), .B(OR4_1266_Y), .C(OR4_1944_Y), .D(
        OR4_2215_Y), .Y(OR4_297_Y));
    OR4 OR4_2270 (.A(\B_DOUT_TEMPR60[8] ), .B(\B_DOUT_TEMPR61[8] ), .C(
        \B_DOUT_TEMPR62[8] ), .D(\B_DOUT_TEMPR63[8] ), .Y(OR4_2270_Y));
    OR4 OR4_2513 (.A(OR4_340_Y), .B(OR4_651_Y), .C(OR4_2231_Y), .D(
        OR4_122_Y), .Y(OR4_2513_Y));
    OR4 OR4_3033 (.A(\A_DOUT_TEMPR32[33] ), .B(\A_DOUT_TEMPR33[33] ), 
        .C(\A_DOUT_TEMPR34[33] ), .D(\A_DOUT_TEMPR35[33] ), .Y(
        OR4_3033_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%72%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R72C6 (
        .A_DOUT({nc12900, nc12901, nc12902, nc12903, nc12904, nc12905, 
        nc12906, nc12907, nc12908, nc12909, nc12910, nc12911, nc12912, 
        nc12913, nc12914, \A_DOUT_TEMPR72[34] , \A_DOUT_TEMPR72[33] , 
        \A_DOUT_TEMPR72[32] , \A_DOUT_TEMPR72[31] , 
        \A_DOUT_TEMPR72[30] }), .B_DOUT({nc12915, nc12916, nc12917, 
        nc12918, nc12919, nc12920, nc12921, nc12922, nc12923, nc12924, 
        nc12925, nc12926, nc12927, nc12928, nc12929, 
        \B_DOUT_TEMPR72[34] , \B_DOUT_TEMPR72[33] , 
        \B_DOUT_TEMPR72[32] , \B_DOUT_TEMPR72[31] , 
        \B_DOUT_TEMPR72[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[72][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2426 (.A(\A_DOUT_TEMPR40[39] ), .B(\A_DOUT_TEMPR41[39] ), 
        .C(\A_DOUT_TEMPR42[39] ), .D(\A_DOUT_TEMPR43[39] ), .Y(
        OR4_2426_Y));
    OR4 OR4_2161 (.A(\B_DOUT_TEMPR4[27] ), .B(\B_DOUT_TEMPR5[27] ), .C(
        \B_DOUT_TEMPR6[27] ), .D(\B_DOUT_TEMPR7[27] ), .Y(OR4_2161_Y));
    OR2 OR2_22 (.A(\A_DOUT_TEMPR72[19] ), .B(\A_DOUT_TEMPR73[19] ), .Y(
        OR2_22_Y));
    OR4 OR4_1327 (.A(\A_DOUT_TEMPR8[2] ), .B(\A_DOUT_TEMPR9[2] ), .C(
        \A_DOUT_TEMPR10[2] ), .D(\A_DOUT_TEMPR11[2] ), .Y(OR4_1327_Y));
    OR4 OR4_1222 (.A(\B_DOUT_TEMPR64[19] ), .B(\B_DOUT_TEMPR65[19] ), 
        .C(\B_DOUT_TEMPR66[19] ), .D(\B_DOUT_TEMPR67[19] ), .Y(
        OR4_1222_Y));
    OR4 OR4_2113 (.A(OR4_613_Y), .B(OR4_2156_Y), .C(OR4_3021_Y), .D(
        OR4_2035_Y), .Y(OR4_2113_Y));
    OR4 OR4_814 (.A(\A_DOUT_TEMPR44[25] ), .B(\A_DOUT_TEMPR45[25] ), 
        .C(\A_DOUT_TEMPR46[25] ), .D(\A_DOUT_TEMPR47[25] ), .Y(
        OR4_814_Y));
    OR4 OR4_1662 (.A(\A_DOUT_TEMPR99[20] ), .B(\A_DOUT_TEMPR100[20] ), 
        .C(\A_DOUT_TEMPR101[20] ), .D(\A_DOUT_TEMPR102[20] ), .Y(
        OR4_1662_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%79%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R79C0 (
        .A_DOUT({nc12930, nc12931, nc12932, nc12933, nc12934, nc12935, 
        nc12936, nc12937, nc12938, nc12939, nc12940, nc12941, nc12942, 
        nc12943, nc12944, \A_DOUT_TEMPR79[4] , \A_DOUT_TEMPR79[3] , 
        \A_DOUT_TEMPR79[2] , \A_DOUT_TEMPR79[1] , \A_DOUT_TEMPR79[0] })
        , .B_DOUT({nc12945, nc12946, nc12947, nc12948, nc12949, 
        nc12950, nc12951, nc12952, nc12953, nc12954, nc12955, nc12956, 
        nc12957, nc12958, nc12959, \B_DOUT_TEMPR79[4] , 
        \B_DOUT_TEMPR79[3] , \B_DOUT_TEMPR79[2] , \B_DOUT_TEMPR79[1] , 
        \B_DOUT_TEMPR79[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[79][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_385 (.A(\B_DOUT_TEMPR24[20] ), .B(\B_DOUT_TEMPR25[20] ), 
        .C(\B_DOUT_TEMPR26[20] ), .D(\B_DOUT_TEMPR27[20] ), .Y(
        OR4_385_Y));
    OR4 OR4_992 (.A(OR4_1772_Y), .B(OR4_61_Y), .C(OR4_2768_Y), .D(
        OR4_755_Y), .Y(OR4_992_Y));
    OR4 OR4_367 (.A(\A_DOUT_TEMPR40[35] ), .B(\A_DOUT_TEMPR41[35] ), 
        .C(\A_DOUT_TEMPR42[35] ), .D(\A_DOUT_TEMPR43[35] ), .Y(
        OR4_367_Y));
    OR4 OR4_512 (.A(\A_DOUT_TEMPR115[35] ), .B(\A_DOUT_TEMPR116[35] ), 
        .C(\A_DOUT_TEMPR117[35] ), .D(\A_DOUT_TEMPR118[35] ), .Y(
        OR4_512_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%91%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R91C7 (
        .A_DOUT({nc12960, nc12961, nc12962, nc12963, nc12964, nc12965, 
        nc12966, nc12967, nc12968, nc12969, nc12970, nc12971, nc12972, 
        nc12973, nc12974, \A_DOUT_TEMPR91[39] , \A_DOUT_TEMPR91[38] , 
        \A_DOUT_TEMPR91[37] , \A_DOUT_TEMPR91[36] , 
        \A_DOUT_TEMPR91[35] }), .B_DOUT({nc12975, nc12976, nc12977, 
        nc12978, nc12979, nc12980, nc12981, nc12982, nc12983, nc12984, 
        nc12985, nc12986, nc12987, nc12988, nc12989, 
        \B_DOUT_TEMPR91[39] , \B_DOUT_TEMPR91[38] , 
        \B_DOUT_TEMPR91[37] , \B_DOUT_TEMPR91[36] , 
        \B_DOUT_TEMPR91[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[91][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2630 (.A(\A_DOUT_TEMPR40[20] ), .B(\A_DOUT_TEMPR41[20] ), 
        .C(\A_DOUT_TEMPR42[20] ), .D(\A_DOUT_TEMPR43[20] ), .Y(
        OR4_2630_Y));
    OR4 OR4_2065 (.A(\A_DOUT_TEMPR16[32] ), .B(\A_DOUT_TEMPR17[32] ), 
        .C(\A_DOUT_TEMPR18[32] ), .D(\A_DOUT_TEMPR19[32] ), .Y(
        OR4_2065_Y));
    OR4 OR4_2012 (.A(\A_DOUT_TEMPR99[4] ), .B(\A_DOUT_TEMPR100[4] ), 
        .C(\A_DOUT_TEMPR101[4] ), .D(\A_DOUT_TEMPR102[4] ), .Y(
        OR4_2012_Y));
    OR4 OR4_195 (.A(\B_DOUT_TEMPR24[37] ), .B(\B_DOUT_TEMPR25[37] ), 
        .C(\B_DOUT_TEMPR26[37] ), .D(\B_DOUT_TEMPR27[37] ), .Y(
        OR4_195_Y));
    OR4 OR4_1118 (.A(\A_DOUT_TEMPR60[20] ), .B(\A_DOUT_TEMPR61[20] ), 
        .C(\A_DOUT_TEMPR62[20] ), .D(\A_DOUT_TEMPR63[20] ), .Y(
        OR4_1118_Y));
    OR4 OR4_1250 (.A(\A_DOUT_TEMPR83[19] ), .B(\A_DOUT_TEMPR84[19] ), 
        .C(\A_DOUT_TEMPR85[19] ), .D(\A_DOUT_TEMPR86[19] ), .Y(
        OR4_1250_Y));
    OR4 OR4_1962 (.A(\B_DOUT_TEMPR12[24] ), .B(\B_DOUT_TEMPR13[24] ), 
        .C(\B_DOUT_TEMPR14[24] ), .D(\B_DOUT_TEMPR15[24] ), .Y(
        OR4_1962_Y));
    OR4 OR4_868 (.A(\A_DOUT_TEMPR28[39] ), .B(\A_DOUT_TEMPR29[39] ), 
        .C(\A_DOUT_TEMPR30[39] ), .D(\A_DOUT_TEMPR31[39] ), .Y(
        OR4_868_Y));
    OR4 OR4_2038 (.A(\B_DOUT_TEMPR4[37] ), .B(\B_DOUT_TEMPR5[37] ), .C(
        \B_DOUT_TEMPR6[37] ), .D(\B_DOUT_TEMPR7[37] ), .Y(OR4_2038_Y));
    OR4 OR4_2376 (.A(\B_DOUT_TEMPR79[13] ), .B(\B_DOUT_TEMPR80[13] ), 
        .C(\B_DOUT_TEMPR81[13] ), .D(\B_DOUT_TEMPR82[13] ), .Y(
        OR4_2376_Y));
    OR4 OR4_661 (.A(OR4_324_Y), .B(OR4_1322_Y), .C(OR4_341_Y), .D(
        OR4_1894_Y), .Y(OR4_661_Y));
    OR4 OR4_1630 (.A(\B_DOUT_TEMPR68[13] ), .B(\B_DOUT_TEMPR69[13] ), 
        .C(\B_DOUT_TEMPR70[13] ), .D(\B_DOUT_TEMPR71[13] ), .Y(
        OR4_1630_Y));
    OR4 OR4_990 (.A(OR4_2607_Y), .B(OR4_1370_Y), .C(OR4_959_Y), .D(
        OR4_2615_Y), .Y(OR4_990_Y));
    OR4 OR4_3018 (.A(\A_DOUT_TEMPR91[24] ), .B(\A_DOUT_TEMPR92[24] ), 
        .C(\A_DOUT_TEMPR93[24] ), .D(\A_DOUT_TEMPR94[24] ), .Y(
        OR4_3018_Y));
    OR4 OR4_2725 (.A(\A_DOUT_TEMPR28[5] ), .B(\A_DOUT_TEMPR29[5] ), .C(
        \A_DOUT_TEMPR30[5] ), .D(\A_DOUT_TEMPR31[5] ), .Y(OR4_2725_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%75%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R75C6 (
        .A_DOUT({nc12990, nc12991, nc12992, nc12993, nc12994, nc12995, 
        nc12996, nc12997, nc12998, nc12999, nc13000, nc13001, nc13002, 
        nc13003, nc13004, \A_DOUT_TEMPR75[34] , \A_DOUT_TEMPR75[33] , 
        \A_DOUT_TEMPR75[32] , \A_DOUT_TEMPR75[31] , 
        \A_DOUT_TEMPR75[30] }), .B_DOUT({nc13005, nc13006, nc13007, 
        nc13008, nc13009, nc13010, nc13011, nc13012, nc13013, nc13014, 
        nc13015, nc13016, nc13017, nc13018, nc13019, 
        \B_DOUT_TEMPR75[34] , \B_DOUT_TEMPR75[33] , 
        \B_DOUT_TEMPR75[32] , \B_DOUT_TEMPR75[31] , 
        \B_DOUT_TEMPR75[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[75][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%85%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R85C0 (
        .A_DOUT({nc13020, nc13021, nc13022, nc13023, nc13024, nc13025, 
        nc13026, nc13027, nc13028, nc13029, nc13030, nc13031, nc13032, 
        nc13033, nc13034, \A_DOUT_TEMPR85[4] , \A_DOUT_TEMPR85[3] , 
        \A_DOUT_TEMPR85[2] , \A_DOUT_TEMPR85[1] , \A_DOUT_TEMPR85[0] })
        , .B_DOUT({nc13035, nc13036, nc13037, nc13038, nc13039, 
        nc13040, nc13041, nc13042, nc13043, nc13044, nc13045, nc13046, 
        nc13047, nc13048, nc13049, \B_DOUT_TEMPR85[4] , 
        \B_DOUT_TEMPR85[3] , \B_DOUT_TEMPR85[2] , \B_DOUT_TEMPR85[1] , 
        \B_DOUT_TEMPR85[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[85][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_477 (.A(\B_DOUT_TEMPR12[6] ), .B(\B_DOUT_TEMPR13[6] ), .C(
        \B_DOUT_TEMPR14[6] ), .D(\B_DOUT_TEMPR15[6] ), .Y(OR4_477_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%56%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R56C1 (
        .A_DOUT({nc13050, nc13051, nc13052, nc13053, nc13054, nc13055, 
        nc13056, nc13057, nc13058, nc13059, nc13060, nc13061, nc13062, 
        nc13063, nc13064, \A_DOUT_TEMPR56[9] , \A_DOUT_TEMPR56[8] , 
        \A_DOUT_TEMPR56[7] , \A_DOUT_TEMPR56[6] , \A_DOUT_TEMPR56[5] })
        , .B_DOUT({nc13065, nc13066, nc13067, nc13068, nc13069, 
        nc13070, nc13071, nc13072, nc13073, nc13074, nc13075, nc13076, 
        nc13077, nc13078, nc13079, \B_DOUT_TEMPR56[9] , 
        \B_DOUT_TEMPR56[8] , \B_DOUT_TEMPR56[7] , \B_DOUT_TEMPR56[6] , 
        \B_DOUT_TEMPR56[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[56][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_223 (.A(\A_DOUT_TEMPR48[30] ), .B(\A_DOUT_TEMPR49[30] ), 
        .C(\A_DOUT_TEMPR50[30] ), .D(\A_DOUT_TEMPR51[30] ), .Y(
        OR4_223_Y));
    OR4 OR4_1038 (.A(OR4_2732_Y), .B(OR4_1668_Y), .C(OR4_2297_Y), .D(
        OR4_1487_Y), .Y(OR4_1038_Y));
    OR4 OR4_1424 (.A(\B_DOUT_TEMPR24[18] ), .B(\B_DOUT_TEMPR25[18] ), 
        .C(\B_DOUT_TEMPR26[18] ), .D(\B_DOUT_TEMPR27[18] ), .Y(
        OR4_1424_Y));
    OR4 OR4_321 (.A(\A_DOUT_TEMPR103[13] ), .B(\A_DOUT_TEMPR104[13] ), 
        .C(\A_DOUT_TEMPR105[13] ), .D(\A_DOUT_TEMPR106[13] ), .Y(
        OR4_321_Y));
    OR4 OR4_825 (.A(\B_DOUT_TEMPR24[38] ), .B(\B_DOUT_TEMPR25[38] ), 
        .C(\B_DOUT_TEMPR26[38] ), .D(\B_DOUT_TEMPR27[38] ), .Y(
        OR4_825_Y));
    OR4 OR4_1813 (.A(\B_DOUT_TEMPR44[23] ), .B(\B_DOUT_TEMPR45[23] ), 
        .C(\B_DOUT_TEMPR46[23] ), .D(\B_DOUT_TEMPR47[23] ), .Y(
        OR4_1813_Y));
    OR4 OR4_46 (.A(\B_DOUT_TEMPR32[7] ), .B(\B_DOUT_TEMPR33[7] ), .C(
        \B_DOUT_TEMPR34[7] ), .D(\B_DOUT_TEMPR35[7] ), .Y(OR4_46_Y));
    OR4 OR4_123 (.A(\B_DOUT_TEMPR20[34] ), .B(\B_DOUT_TEMPR21[34] ), 
        .C(\B_DOUT_TEMPR22[34] ), .D(\B_DOUT_TEMPR23[34] ), .Y(
        OR4_123_Y));
    OR4 OR4_439 (.A(OR4_593_Y), .B(OR4_2980_Y), .C(OR4_2484_Y), .D(
        OR4_2806_Y), .Y(OR4_439_Y));
    OR4 OR4_3031 (.A(\B_DOUT_TEMPR83[23] ), .B(\B_DOUT_TEMPR84[23] ), 
        .C(\B_DOUT_TEMPR85[23] ), .D(\B_DOUT_TEMPR86[23] ), .Y(
        OR4_3031_Y));
    OR4 OR4_2867 (.A(OR4_3_Y), .B(OR4_1329_Y), .C(OR4_978_Y), .D(
        OR4_2012_Y), .Y(OR4_2867_Y));
    OR4 OR4_464 (.A(\B_DOUT_TEMPR36[19] ), .B(\B_DOUT_TEMPR37[19] ), 
        .C(\B_DOUT_TEMPR38[19] ), .D(\B_DOUT_TEMPR39[19] ), .Y(
        OR4_464_Y));
    OR4 OR4_1356 (.A(\B_DOUT_TEMPR4[31] ), .B(\B_DOUT_TEMPR5[31] ), .C(
        \B_DOUT_TEMPR6[31] ), .D(\B_DOUT_TEMPR7[31] ), .Y(OR4_1356_Y));
    OR4 OR4_2901 (.A(OR4_2571_Y), .B(OR4_1574_Y), .C(OR4_2524_Y), .D(
        OR4_701_Y), .Y(OR4_2901_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%56%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R56C2 (
        .A_DOUT({nc13080, nc13081, nc13082, nc13083, nc13084, nc13085, 
        nc13086, nc13087, nc13088, nc13089, nc13090, nc13091, nc13092, 
        nc13093, nc13094, \A_DOUT_TEMPR56[14] , \A_DOUT_TEMPR56[13] , 
        \A_DOUT_TEMPR56[12] , \A_DOUT_TEMPR56[11] , 
        \A_DOUT_TEMPR56[10] }), .B_DOUT({nc13095, nc13096, nc13097, 
        nc13098, nc13099, nc13100, nc13101, nc13102, nc13103, nc13104, 
        nc13105, nc13106, nc13107, nc13108, nc13109, 
        \B_DOUT_TEMPR56[14] , \B_DOUT_TEMPR56[13] , 
        \B_DOUT_TEMPR56[12] , \B_DOUT_TEMPR56[11] , 
        \B_DOUT_TEMPR56[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[56][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1719 (.A(\B_DOUT_TEMPR79[20] ), .B(\B_DOUT_TEMPR80[20] ), 
        .C(\B_DOUT_TEMPR81[20] ), .D(\B_DOUT_TEMPR82[20] ), .Y(
        OR4_1719_Y));
    OR4 OR4_1695 (.A(OR4_389_Y), .B(OR4_770_Y), .C(OR4_1519_Y), .D(
        OR4_2321_Y), .Y(OR4_1695_Y));
    OR4 OR4_2158 (.A(OR4_143_Y), .B(OR4_3016_Y), .C(OR4_835_Y), .D(
        OR4_2026_Y), .Y(OR4_2158_Y));
    OR4 OR4_2044 (.A(\B_DOUT_TEMPR103[35] ), .B(\B_DOUT_TEMPR104[35] ), 
        .C(\B_DOUT_TEMPR105[35] ), .D(\B_DOUT_TEMPR106[35] ), .Y(
        OR4_2044_Y));
    OR4 OR4_880 (.A(\B_DOUT_TEMPR56[9] ), .B(\B_DOUT_TEMPR57[9] ), .C(
        \B_DOUT_TEMPR58[9] ), .D(\B_DOUT_TEMPR59[9] ), .Y(OR4_880_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%50%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R50C6 (
        .A_DOUT({nc13110, nc13111, nc13112, nc13113, nc13114, nc13115, 
        nc13116, nc13117, nc13118, nc13119, nc13120, nc13121, nc13122, 
        nc13123, nc13124, \A_DOUT_TEMPR50[34] , \A_DOUT_TEMPR50[33] , 
        \A_DOUT_TEMPR50[32] , \A_DOUT_TEMPR50[31] , 
        \A_DOUT_TEMPR50[30] }), .B_DOUT({nc13125, nc13126, nc13127, 
        nc13128, nc13129, nc13130, nc13131, nc13132, nc13133, nc13134, 
        nc13135, nc13136, nc13137, nc13138, nc13139, 
        \B_DOUT_TEMPR50[34] , \B_DOUT_TEMPR50[33] , 
        \B_DOUT_TEMPR50[32] , \B_DOUT_TEMPR50[31] , 
        \B_DOUT_TEMPR50[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2046 (.A(\B_DOUT_TEMPR60[32] ), .B(\B_DOUT_TEMPR61[32] ), 
        .C(\B_DOUT_TEMPR62[32] ), .D(\B_DOUT_TEMPR63[32] ), .Y(
        OR4_2046_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%24%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R24C0 (
        .A_DOUT({nc13140, nc13141, nc13142, nc13143, nc13144, nc13145, 
        nc13146, nc13147, nc13148, nc13149, nc13150, nc13151, nc13152, 
        nc13153, nc13154, \A_DOUT_TEMPR24[4] , \A_DOUT_TEMPR24[3] , 
        \A_DOUT_TEMPR24[2] , \A_DOUT_TEMPR24[1] , \A_DOUT_TEMPR24[0] })
        , .B_DOUT({nc13155, nc13156, nc13157, nc13158, nc13159, 
        nc13160, nc13161, nc13162, nc13163, nc13164, nc13165, nc13166, 
        nc13167, nc13168, nc13169, \B_DOUT_TEMPR24[4] , 
        \B_DOUT_TEMPR24[3] , \B_DOUT_TEMPR24[2] , \B_DOUT_TEMPR24[1] , 
        \B_DOUT_TEMPR24[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%50%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R50C5 (
        .A_DOUT({nc13170, nc13171, nc13172, nc13173, nc13174, nc13175, 
        nc13176, nc13177, nc13178, nc13179, nc13180, nc13181, nc13182, 
        nc13183, nc13184, \A_DOUT_TEMPR50[29] , \A_DOUT_TEMPR50[28] , 
        \A_DOUT_TEMPR50[27] , \A_DOUT_TEMPR50[26] , 
        \A_DOUT_TEMPR50[25] }), .B_DOUT({nc13185, nc13186, nc13187, 
        nc13188, nc13189, nc13190, nc13191, nc13192, nc13193, nc13194, 
        nc13195, nc13196, nc13197, nc13198, nc13199, 
        \B_DOUT_TEMPR50[29] , \B_DOUT_TEMPR50[28] , 
        \B_DOUT_TEMPR50[27] , \B_DOUT_TEMPR50[26] , 
        \B_DOUT_TEMPR50[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_580 (.A(OR4_2448_Y), .B(OR4_1471_Y), .C(OR4_1673_Y), .D(
        OR4_1485_Y), .Y(OR4_580_Y));
    OR4 OR4_1116 (.A(\B_DOUT_TEMPR75[20] ), .B(\B_DOUT_TEMPR76[20] ), 
        .C(\B_DOUT_TEMPR77[20] ), .D(\B_DOUT_TEMPR78[20] ), .Y(
        OR4_1116_Y));
    OR4 OR4_2192 (.A(\B_DOUT_TEMPR24[27] ), .B(\B_DOUT_TEMPR25[27] ), 
        .C(\B_DOUT_TEMPR26[27] ), .D(\B_DOUT_TEMPR27[27] ), .Y(
        OR4_2192_Y));
    OR4 OR4_2134 (.A(\B_DOUT_TEMPR115[15] ), .B(\B_DOUT_TEMPR116[15] ), 
        .C(\B_DOUT_TEMPR117[15] ), .D(\B_DOUT_TEMPR118[15] ), .Y(
        OR4_2134_Y));
    OR4 OR4_1518 (.A(OR4_2388_Y), .B(OR4_335_Y), .C(OR4_1051_Y), .D(
        OR4_2710_Y), .Y(OR4_1518_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%107%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R107C5 (
        .A_DOUT({nc13200, nc13201, nc13202, nc13203, nc13204, nc13205, 
        nc13206, nc13207, nc13208, nc13209, nc13210, nc13211, nc13212, 
        nc13213, nc13214, \A_DOUT_TEMPR107[29] , \A_DOUT_TEMPR107[28] , 
        \A_DOUT_TEMPR107[27] , \A_DOUT_TEMPR107[26] , 
        \A_DOUT_TEMPR107[25] }), .B_DOUT({nc13215, nc13216, nc13217, 
        nc13218, nc13219, nc13220, nc13221, nc13222, nc13223, nc13224, 
        nc13225, nc13226, nc13227, nc13228, nc13229, 
        \B_DOUT_TEMPR107[29] , \B_DOUT_TEMPR107[28] , 
        \B_DOUT_TEMPR107[27] , \B_DOUT_TEMPR107[26] , 
        \B_DOUT_TEMPR107[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[107][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_24 (.A(\A_DOUT_TEMPR72[25] ), .B(\A_DOUT_TEMPR73[25] ), .Y(
        OR2_24_Y));
    OR4 OR4_131 (.A(OR4_2174_Y), .B(OR4_2733_Y), .C(OR4_2264_Y), .D(
        OR4_946_Y), .Y(OR4_131_Y));
    OR4 OR4_2853 (.A(\B_DOUT_TEMPR103[5] ), .B(\B_DOUT_TEMPR104[5] ), 
        .C(\B_DOUT_TEMPR105[5] ), .D(\B_DOUT_TEMPR106[5] ), .Y(
        OR4_2853_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_21 (.A(B_BLK_EN), .B(B_ADDR[18]), .C(
        B_ADDR[17]), .Y(CFG3_21_Y));
    OR4 OR4_722 (.A(\A_DOUT_TEMPR52[33] ), .B(\A_DOUT_TEMPR53[33] ), 
        .C(\A_DOUT_TEMPR54[33] ), .D(\A_DOUT_TEMPR55[33] ), .Y(
        OR4_722_Y));
    OR4 OR4_1586 (.A(\A_DOUT_TEMPR111[4] ), .B(\A_DOUT_TEMPR112[4] ), 
        .C(\A_DOUT_TEMPR113[4] ), .D(\A_DOUT_TEMPR114[4] ), .Y(
        OR4_1586_Y));
    OR4 OR4_784 (.A(\B_DOUT_TEMPR79[23] ), .B(\B_DOUT_TEMPR80[23] ), 
        .C(\B_DOUT_TEMPR81[23] ), .D(\B_DOUT_TEMPR82[23] ), .Y(
        OR4_784_Y));
    OR4 OR4_2343 (.A(\A_DOUT_TEMPR12[22] ), .B(\A_DOUT_TEMPR13[22] ), 
        .C(\A_DOUT_TEMPR14[22] ), .D(\A_DOUT_TEMPR15[22] ), .Y(
        OR4_2343_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%26%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R26C7 (
        .A_DOUT({nc13230, nc13231, nc13232, nc13233, nc13234, nc13235, 
        nc13236, nc13237, nc13238, nc13239, nc13240, nc13241, nc13242, 
        nc13243, nc13244, \A_DOUT_TEMPR26[39] , \A_DOUT_TEMPR26[38] , 
        \A_DOUT_TEMPR26[37] , \A_DOUT_TEMPR26[36] , 
        \A_DOUT_TEMPR26[35] }), .B_DOUT({nc13245, nc13246, nc13247, 
        nc13248, nc13249, nc13250, nc13251, nc13252, nc13253, nc13254, 
        nc13255, nc13256, nc13257, nc13258, nc13259, 
        \B_DOUT_TEMPR26[39] , \B_DOUT_TEMPR26[38] , 
        \B_DOUT_TEMPR26[37] , \B_DOUT_TEMPR26[36] , 
        \B_DOUT_TEMPR26[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1697 (.A(\A_DOUT_TEMPR24[12] ), .B(\A_DOUT_TEMPR25[12] ), 
        .C(\A_DOUT_TEMPR26[12] ), .D(\A_DOUT_TEMPR27[12] ), .Y(
        OR4_1697_Y));
    OR4 OR4_326 (.A(\A_DOUT_TEMPR103[29] ), .B(\A_DOUT_TEMPR104[29] ), 
        .C(\A_DOUT_TEMPR105[29] ), .D(\A_DOUT_TEMPR106[29] ), .Y(
        OR4_326_Y));
    OR4 OR4_1787 (.A(\B_DOUT_TEMPR103[7] ), .B(\B_DOUT_TEMPR104[7] ), 
        .C(\B_DOUT_TEMPR105[7] ), .D(\B_DOUT_TEMPR106[7] ), .Y(
        OR4_1787_Y));
    OR4 OR4_407 (.A(\B_DOUT_TEMPR32[32] ), .B(\B_DOUT_TEMPR33[32] ), 
        .C(\B_DOUT_TEMPR34[32] ), .D(\B_DOUT_TEMPR35[32] ), .Y(
        OR4_407_Y));
    OR4 OR4_1134 (.A(\B_DOUT_TEMPR20[5] ), .B(\B_DOUT_TEMPR21[5] ), .C(
        \B_DOUT_TEMPR22[5] ), .D(\B_DOUT_TEMPR23[5] ), .Y(OR4_1134_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%42%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R42C5 (
        .A_DOUT({nc13260, nc13261, nc13262, nc13263, nc13264, nc13265, 
        nc13266, nc13267, nc13268, nc13269, nc13270, nc13271, nc13272, 
        nc13273, nc13274, \A_DOUT_TEMPR42[29] , \A_DOUT_TEMPR42[28] , 
        \A_DOUT_TEMPR42[27] , \A_DOUT_TEMPR42[26] , 
        \A_DOUT_TEMPR42[25] }), .B_DOUT({nc13275, nc13276, nc13277, 
        nc13278, nc13279, nc13280, nc13281, nc13282, nc13283, nc13284, 
        nc13285, nc13286, nc13287, nc13288, nc13289, 
        \B_DOUT_TEMPR42[29] , \B_DOUT_TEMPR42[28] , 
        \B_DOUT_TEMPR42[27] , \B_DOUT_TEMPR42[26] , 
        \B_DOUT_TEMPR42[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[42][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1581 (.A(\B_DOUT_TEMPR12[16] ), .B(\B_DOUT_TEMPR13[16] ), 
        .C(\B_DOUT_TEMPR14[16] ), .D(\B_DOUT_TEMPR15[16] ), .Y(
        OR4_1581_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%89%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R89C1 (
        .A_DOUT({nc13290, nc13291, nc13292, nc13293, nc13294, nc13295, 
        nc13296, nc13297, nc13298, nc13299, nc13300, nc13301, nc13302, 
        nc13303, nc13304, \A_DOUT_TEMPR89[9] , \A_DOUT_TEMPR89[8] , 
        \A_DOUT_TEMPR89[7] , \A_DOUT_TEMPR89[6] , \A_DOUT_TEMPR89[5] })
        , .B_DOUT({nc13305, nc13306, nc13307, nc13308, nc13309, 
        nc13310, nc13311, nc13312, nc13313, nc13314, nc13315, nc13316, 
        nc13317, nc13318, nc13319, \B_DOUT_TEMPR89[9] , 
        \B_DOUT_TEMPR89[8] , \B_DOUT_TEMPR89[7] , \B_DOUT_TEMPR89[6] , 
        \B_DOUT_TEMPR89[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[89][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2759 (.A(\A_DOUT_TEMPR44[7] ), .B(\A_DOUT_TEMPR45[7] ), .C(
        \A_DOUT_TEMPR46[7] ), .D(\A_DOUT_TEMPR47[7] ), .Y(OR4_2759_Y));
    OR4 OR4_2472 (.A(\B_DOUT_TEMPR107[28] ), .B(\B_DOUT_TEMPR108[28] ), 
        .C(\B_DOUT_TEMPR109[28] ), .D(\B_DOUT_TEMPR110[28] ), .Y(
        OR4_2472_Y));
    OR4 OR4_2203 (.A(OR4_2444_Y), .B(OR4_845_Y), .C(OR2_8_Y), .D(
        \A_DOUT_TEMPR74[8] ), .Y(OR4_2203_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%27%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R27C6 (
        .A_DOUT({nc13320, nc13321, nc13322, nc13323, nc13324, nc13325, 
        nc13326, nc13327, nc13328, nc13329, nc13330, nc13331, nc13332, 
        nc13333, nc13334, \A_DOUT_TEMPR27[34] , \A_DOUT_TEMPR27[33] , 
        \A_DOUT_TEMPR27[32] , \A_DOUT_TEMPR27[31] , 
        \A_DOUT_TEMPR27[30] }), .B_DOUT({nc13335, nc13336, nc13337, 
        nc13338, nc13339, nc13340, nc13341, nc13342, nc13343, nc13344, 
        nc13345, nc13346, nc13347, nc13348, nc13349, 
        \B_DOUT_TEMPR27[34] , \B_DOUT_TEMPR27[33] , 
        \B_DOUT_TEMPR27[32] , \B_DOUT_TEMPR27[31] , 
        \B_DOUT_TEMPR27[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2478 (.A(\A_DOUT_TEMPR64[15] ), .B(\A_DOUT_TEMPR65[15] ), 
        .C(\A_DOUT_TEMPR66[15] ), .D(\A_DOUT_TEMPR67[15] ), .Y(
        OR4_2478_Y));
    OR4 OR4_1469 (.A(OR4_9_Y), .B(OR4_1589_Y), .C(OR4_2809_Y), .D(
        OR4_2506_Y), .Y(OR4_1469_Y));
    OR4 OR4_527 (.A(\B_DOUT_TEMPR4[12] ), .B(\B_DOUT_TEMPR5[12] ), .C(
        \B_DOUT_TEMPR6[12] ), .D(\B_DOUT_TEMPR7[12] ), .Y(OR4_527_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%36%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R36C1 (
        .A_DOUT({nc13350, nc13351, nc13352, nc13353, nc13354, nc13355, 
        nc13356, nc13357, nc13358, nc13359, nc13360, nc13361, nc13362, 
        nc13363, nc13364, \A_DOUT_TEMPR36[9] , \A_DOUT_TEMPR36[8] , 
        \A_DOUT_TEMPR36[7] , \A_DOUT_TEMPR36[6] , \A_DOUT_TEMPR36[5] })
        , .B_DOUT({nc13365, nc13366, nc13367, nc13368, nc13369, 
        nc13370, nc13371, nc13372, nc13373, nc13374, nc13375, nc13376, 
        nc13377, nc13378, nc13379, \B_DOUT_TEMPR36[9] , 
        \B_DOUT_TEMPR36[8] , \B_DOUT_TEMPR36[7] , \B_DOUT_TEMPR36[6] , 
        \B_DOUT_TEMPR36[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%97%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R97C0 (
        .A_DOUT({nc13380, nc13381, nc13382, nc13383, nc13384, nc13385, 
        nc13386, nc13387, nc13388, nc13389, nc13390, nc13391, nc13392, 
        nc13393, nc13394, \A_DOUT_TEMPR97[4] , \A_DOUT_TEMPR97[3] , 
        \A_DOUT_TEMPR97[2] , \A_DOUT_TEMPR97[1] , \A_DOUT_TEMPR97[0] })
        , .B_DOUT({nc13395, nc13396, nc13397, nc13398, nc13399, 
        nc13400, nc13401, nc13402, nc13403, nc13404, nc13405, nc13406, 
        nc13407, nc13408, nc13409, \B_DOUT_TEMPR97[4] , 
        \B_DOUT_TEMPR97[3] , \B_DOUT_TEMPR97[2] , \B_DOUT_TEMPR97[1] , 
        \B_DOUT_TEMPR97[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[97][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%42%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R42C1 (
        .A_DOUT({nc13410, nc13411, nc13412, nc13413, nc13414, nc13415, 
        nc13416, nc13417, nc13418, nc13419, nc13420, nc13421, nc13422, 
        nc13423, nc13424, \A_DOUT_TEMPR42[9] , \A_DOUT_TEMPR42[8] , 
        \A_DOUT_TEMPR42[7] , \A_DOUT_TEMPR42[6] , \A_DOUT_TEMPR42[5] })
        , .B_DOUT({nc13425, nc13426, nc13427, nc13428, nc13429, 
        nc13430, nc13431, nc13432, nc13433, nc13434, nc13435, nc13436, 
        nc13437, nc13438, nc13439, \B_DOUT_TEMPR42[9] , 
        \B_DOUT_TEMPR42[8] , \B_DOUT_TEMPR42[7] , \B_DOUT_TEMPR42[6] , 
        \B_DOUT_TEMPR42[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[42][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%19%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R19C7 (
        .A_DOUT({nc13440, nc13441, nc13442, nc13443, nc13444, nc13445, 
        nc13446, nc13447, nc13448, nc13449, nc13450, nc13451, nc13452, 
        nc13453, nc13454, \A_DOUT_TEMPR19[39] , \A_DOUT_TEMPR19[38] , 
        \A_DOUT_TEMPR19[37] , \A_DOUT_TEMPR19[36] , 
        \A_DOUT_TEMPR19[35] }), .B_DOUT({nc13455, nc13456, nc13457, 
        nc13458, nc13459, nc13460, nc13461, nc13462, nc13463, nc13464, 
        nc13465, nc13466, nc13467, nc13468, nc13469, 
        \B_DOUT_TEMPR19[39] , \B_DOUT_TEMPR19[38] , 
        \B_DOUT_TEMPR19[37] , \B_DOUT_TEMPR19[36] , 
        \B_DOUT_TEMPR19[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_243 (.A(\B_DOUT_TEMPR99[6] ), .B(\B_DOUT_TEMPR100[6] ), .C(
        \B_DOUT_TEMPR101[6] ), .D(\B_DOUT_TEMPR102[6] ), .Y(OR4_243_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%112%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R112C2 (
        .A_DOUT({nc13470, nc13471, nc13472, nc13473, nc13474, nc13475, 
        nc13476, nc13477, nc13478, nc13479, nc13480, nc13481, nc13482, 
        nc13483, nc13484, \A_DOUT_TEMPR112[14] , \A_DOUT_TEMPR112[13] , 
        \A_DOUT_TEMPR112[12] , \A_DOUT_TEMPR112[11] , 
        \A_DOUT_TEMPR112[10] }), .B_DOUT({nc13485, nc13486, nc13487, 
        nc13488, nc13489, nc13490, nc13491, nc13492, nc13493, nc13494, 
        nc13495, nc13496, nc13497, nc13498, nc13499, 
        \B_DOUT_TEMPR112[14] , \B_DOUT_TEMPR112[13] , 
        \B_DOUT_TEMPR112[12] , \B_DOUT_TEMPR112[11] , 
        \B_DOUT_TEMPR112[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[112][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1224 (.A(\B_DOUT_TEMPR56[27] ), .B(\B_DOUT_TEMPR57[27] ), 
        .C(\B_DOUT_TEMPR58[27] ), .D(\B_DOUT_TEMPR59[27] ), .Y(
        OR4_1224_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%6%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R6C6 (
        .A_DOUT({nc13500, nc13501, nc13502, nc13503, nc13504, nc13505, 
        nc13506, nc13507, nc13508, nc13509, nc13510, nc13511, nc13512, 
        nc13513, nc13514, \A_DOUT_TEMPR6[34] , \A_DOUT_TEMPR6[33] , 
        \A_DOUT_TEMPR6[32] , \A_DOUT_TEMPR6[31] , \A_DOUT_TEMPR6[30] })
        , .B_DOUT({nc13515, nc13516, nc13517, nc13518, nc13519, 
        nc13520, nc13521, nc13522, nc13523, nc13524, nc13525, nc13526, 
        nc13527, nc13528, nc13529, \B_DOUT_TEMPR6[34] , 
        \B_DOUT_TEMPR6[33] , \B_DOUT_TEMPR6[32] , \B_DOUT_TEMPR6[31] , 
        \B_DOUT_TEMPR6[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2182 (.A(OR4_2918_Y), .B(OR4_221_Y), .C(OR4_2899_Y), .D(
        OR4_855_Y), .Y(OR4_2182_Y));
    OR4 OR4_341 (.A(OR4_874_Y), .B(OR4_2916_Y), .C(OR4_546_Y), .D(
        OR4_853_Y), .Y(OR4_341_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%89%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R89C2 (
        .A_DOUT({nc13530, nc13531, nc13532, nc13533, nc13534, nc13535, 
        nc13536, nc13537, nc13538, nc13539, nc13540, nc13541, nc13542, 
        nc13543, nc13544, \A_DOUT_TEMPR89[14] , \A_DOUT_TEMPR89[13] , 
        \A_DOUT_TEMPR89[12] , \A_DOUT_TEMPR89[11] , 
        \A_DOUT_TEMPR89[10] }), .B_DOUT({nc13545, nc13546, nc13547, 
        nc13548, nc13549, nc13550, nc13551, nc13552, nc13553, nc13554, 
        nc13555, nc13556, nc13557, nc13558, nc13559, 
        \B_DOUT_TEMPR89[14] , \B_DOUT_TEMPR89[13] , 
        \B_DOUT_TEMPR89[12] , \B_DOUT_TEMPR89[11] , 
        \B_DOUT_TEMPR89[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[89][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_987 (.A(\A_DOUT_TEMPR107[7] ), .B(\A_DOUT_TEMPR108[7] ), 
        .C(\A_DOUT_TEMPR109[7] ), .D(\A_DOUT_TEMPR110[7] ), .Y(
        OR4_987_Y));
    OR4 OR4_2156 (.A(\A_DOUT_TEMPR4[18] ), .B(\A_DOUT_TEMPR5[18] ), .C(
        \A_DOUT_TEMPR6[18] ), .D(\A_DOUT_TEMPR7[18] ), .Y(OR4_2156_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%85%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R85C1 (
        .A_DOUT({nc13560, nc13561, nc13562, nc13563, nc13564, nc13565, 
        nc13566, nc13567, nc13568, nc13569, nc13570, nc13571, nc13572, 
        nc13573, nc13574, \A_DOUT_TEMPR85[9] , \A_DOUT_TEMPR85[8] , 
        \A_DOUT_TEMPR85[7] , \A_DOUT_TEMPR85[6] , \A_DOUT_TEMPR85[5] })
        , .B_DOUT({nc13575, nc13576, nc13577, nc13578, nc13579, 
        nc13580, nc13581, nc13582, nc13583, nc13584, nc13585, nc13586, 
        nc13587, nc13588, nc13589, \B_DOUT_TEMPR85[9] , 
        \B_DOUT_TEMPR85[8] , \B_DOUT_TEMPR85[7] , \B_DOUT_TEMPR85[6] , 
        \B_DOUT_TEMPR85[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[85][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%108%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R108C5 (
        .A_DOUT({nc13590, nc13591, nc13592, nc13593, nc13594, nc13595, 
        nc13596, nc13597, nc13598, nc13599, nc13600, nc13601, nc13602, 
        nc13603, nc13604, \A_DOUT_TEMPR108[29] , \A_DOUT_TEMPR108[28] , 
        \A_DOUT_TEMPR108[27] , \A_DOUT_TEMPR108[26] , 
        \A_DOUT_TEMPR108[25] }), .B_DOUT({nc13605, nc13606, nc13607, 
        nc13608, nc13609, nc13610, nc13611, nc13612, nc13613, nc13614, 
        nc13615, nc13616, nc13617, nc13618, nc13619, 
        \B_DOUT_TEMPR108[29] , \B_DOUT_TEMPR108[28] , 
        \B_DOUT_TEMPR108[27] , \B_DOUT_TEMPR108[26] , 
        \B_DOUT_TEMPR108[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[108][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_845 (.A(\A_DOUT_TEMPR68[8] ), .B(\A_DOUT_TEMPR69[8] ), .C(
        \A_DOUT_TEMPR70[8] ), .D(\A_DOUT_TEMPR71[8] ), .Y(OR4_845_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%8%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R8C4 (
        .A_DOUT({nc13620, nc13621, nc13622, nc13623, nc13624, nc13625, 
        nc13626, nc13627, nc13628, nc13629, nc13630, nc13631, nc13632, 
        nc13633, nc13634, \A_DOUT_TEMPR8[24] , \A_DOUT_TEMPR8[23] , 
        \A_DOUT_TEMPR8[22] , \A_DOUT_TEMPR8[21] , \A_DOUT_TEMPR8[20] })
        , .B_DOUT({nc13635, nc13636, nc13637, nc13638, nc13639, 
        nc13640, nc13641, nc13642, nc13643, nc13644, nc13645, nc13646, 
        nc13647, nc13648, nc13649, \B_DOUT_TEMPR8[24] , 
        \B_DOUT_TEMPR8[23] , \B_DOUT_TEMPR8[22] , \B_DOUT_TEMPR8[21] , 
        \B_DOUT_TEMPR8[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%22%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R22C4 (
        .A_DOUT({nc13650, nc13651, nc13652, nc13653, nc13654, nc13655, 
        nc13656, nc13657, nc13658, nc13659, nc13660, nc13661, nc13662, 
        nc13663, nc13664, \A_DOUT_TEMPR22[24] , \A_DOUT_TEMPR22[23] , 
        \A_DOUT_TEMPR22[22] , \A_DOUT_TEMPR22[21] , 
        \A_DOUT_TEMPR22[20] }), .B_DOUT({nc13665, nc13666, nc13667, 
        nc13668, nc13669, nc13670, nc13671, nc13672, nc13673, nc13674, 
        nc13675, nc13676, nc13677, nc13678, nc13679, 
        \B_DOUT_TEMPR22[24] , \B_DOUT_TEMPR22[23] , 
        \B_DOUT_TEMPR22[22] , \B_DOUT_TEMPR22[21] , 
        \B_DOUT_TEMPR22[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_143 (.A(\A_DOUT_TEMPR16[13] ), .B(\A_DOUT_TEMPR17[13] ), 
        .C(\A_DOUT_TEMPR18[13] ), .D(\A_DOUT_TEMPR19[13] ), .Y(
        OR4_143_Y));
    OR4 OR4_2558 (.A(\B_DOUT_TEMPR83[18] ), .B(\B_DOUT_TEMPR84[18] ), 
        .C(\B_DOUT_TEMPR85[18] ), .D(\B_DOUT_TEMPR86[18] ), .Y(
        OR4_2558_Y));
    OR4 OR4_2835 (.A(OR4_1388_Y), .B(OR4_2258_Y), .C(OR4_4_Y), .D(
        OR4_1518_Y), .Y(OR4_2835_Y));
    OR4 OR4_235 (.A(\B_DOUT_TEMPR36[20] ), .B(\B_DOUT_TEMPR37[20] ), 
        .C(\B_DOUT_TEMPR38[20] ), .D(\B_DOUT_TEMPR39[20] ), .Y(
        OR4_235_Y));
    OR4 OR4_1452 (.A(\A_DOUT_TEMPR60[18] ), .B(\A_DOUT_TEMPR61[18] ), 
        .C(\A_DOUT_TEMPR62[18] ), .D(\A_DOUT_TEMPR63[18] ), .Y(
        OR4_1452_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[8]  (.A(CFG3_11_Y), .B(
        CFG3_15_Y), .Y(\BLKY2[8] ));
    OR4 OR4_1148 (.A(OR4_1461_Y), .B(OR4_2920_Y), .C(OR2_58_Y), .D(
        \A_DOUT_TEMPR74[4] ), .Y(OR4_1148_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%36%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R36C2 (
        .A_DOUT({nc13680, nc13681, nc13682, nc13683, nc13684, nc13685, 
        nc13686, nc13687, nc13688, nc13689, nc13690, nc13691, nc13692, 
        nc13693, nc13694, \A_DOUT_TEMPR36[14] , \A_DOUT_TEMPR36[13] , 
        \A_DOUT_TEMPR36[12] , \A_DOUT_TEMPR36[11] , 
        \A_DOUT_TEMPR36[10] }), .B_DOUT({nc13695, nc13696, nc13697, 
        nc13698, nc13699, nc13700, nc13701, nc13702, nc13703, nc13704, 
        nc13705, nc13706, nc13707, nc13708, nc13709, 
        \B_DOUT_TEMPR36[14] , \B_DOUT_TEMPR36[13] , 
        \B_DOUT_TEMPR36[12] , \B_DOUT_TEMPR36[11] , 
        \B_DOUT_TEMPR36[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENB[8]  (.A(B_WBYTE_EN[4]), .B(
        B_WEN), .Y(\WBYTEENB[8] ));
    OR4 OR4_1835 (.A(\B_DOUT_TEMPR60[24] ), .B(\B_DOUT_TEMPR61[24] ), 
        .C(\B_DOUT_TEMPR62[24] ), .D(\B_DOUT_TEMPR63[24] ), .Y(
        OR4_1835_Y));
    OR4 OR4_1458 (.A(OR4_339_Y), .B(OR4_2741_Y), .C(OR4_1593_Y), .D(
        OR4_2581_Y), .Y(OR4_1458_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%30%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R30C6 (
        .A_DOUT({nc13710, nc13711, nc13712, nc13713, nc13714, nc13715, 
        nc13716, nc13717, nc13718, nc13719, nc13720, nc13721, nc13722, 
        nc13723, nc13724, \A_DOUT_TEMPR30[34] , \A_DOUT_TEMPR30[33] , 
        \A_DOUT_TEMPR30[32] , \A_DOUT_TEMPR30[31] , 
        \A_DOUT_TEMPR30[30] }), .B_DOUT({nc13725, nc13726, nc13727, 
        nc13728, nc13729, nc13730, nc13731, nc13732, nc13733, nc13734, 
        nc13735, nc13736, nc13737, nc13738, nc13739, 
        \B_DOUT_TEMPR30[34] , \B_DOUT_TEMPR30[33] , 
        \B_DOUT_TEMPR30[32] , \B_DOUT_TEMPR30[31] , 
        \B_DOUT_TEMPR30[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2570 (.A(\B_DOUT_TEMPR79[5] ), .B(\B_DOUT_TEMPR80[5] ), .C(
        \B_DOUT_TEMPR81[5] ), .D(\B_DOUT_TEMPR82[5] ), .Y(OR4_2570_Y));
    OR4 OR4_1023 (.A(\B_DOUT_TEMPR36[10] ), .B(\B_DOUT_TEMPR37[10] ), 
        .C(\B_DOUT_TEMPR38[10] ), .D(\B_DOUT_TEMPR39[10] ), .Y(
        OR4_1023_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%30%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R30C5 (
        .A_DOUT({nc13740, nc13741, nc13742, nc13743, nc13744, nc13745, 
        nc13746, nc13747, nc13748, nc13749, nc13750, nc13751, nc13752, 
        nc13753, nc13754, \A_DOUT_TEMPR30[29] , \A_DOUT_TEMPR30[28] , 
        \A_DOUT_TEMPR30[27] , \A_DOUT_TEMPR30[26] , 
        \A_DOUT_TEMPR30[25] }), .B_DOUT({nc13755, nc13756, nc13757, 
        nc13758, nc13759, nc13760, nc13761, nc13762, nc13763, nc13764, 
        nc13765, nc13766, nc13767, nc13768, nc13769, 
        \B_DOUT_TEMPR30[29] , \B_DOUT_TEMPR30[28] , 
        \B_DOUT_TEMPR30[27] , \B_DOUT_TEMPR30[26] , 
        \B_DOUT_TEMPR30[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2526 (.A(OR4_1556_Y), .B(OR4_583_Y), .C(OR4_781_Y), .D(
        OR4_595_Y), .Y(OR4_2526_Y));
    OR4 OR4_586 (.A(\B_DOUT_TEMPR0[15] ), .B(\B_DOUT_TEMPR1[15] ), .C(
        \B_DOUT_TEMPR2[15] ), .D(\B_DOUT_TEMPR3[15] ), .Y(OR4_586_Y));
    OR4 OR4_1360 (.A(OR4_2447_Y), .B(OR4_2247_Y), .C(OR2_51_Y), .D(
        \A_DOUT_TEMPR74[33] ), .Y(OR4_1360_Y));
    OR4 OR4_1467 (.A(\B_DOUT_TEMPR56[29] ), .B(\B_DOUT_TEMPR57[29] ), 
        .C(\B_DOUT_TEMPR58[29] ), .D(\B_DOUT_TEMPR59[29] ), .Y(
        OR4_1467_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%5%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R5C4 (
        .A_DOUT({nc13770, nc13771, nc13772, nc13773, nc13774, nc13775, 
        nc13776, nc13777, nc13778, nc13779, nc13780, nc13781, nc13782, 
        nc13783, nc13784, \A_DOUT_TEMPR5[24] , \A_DOUT_TEMPR5[23] , 
        \A_DOUT_TEMPR5[22] , \A_DOUT_TEMPR5[21] , \A_DOUT_TEMPR5[20] })
        , .B_DOUT({nc13785, nc13786, nc13787, nc13788, nc13789, 
        nc13790, nc13791, nc13792, nc13793, nc13794, nc13795, nc13796, 
        nc13797, nc13798, nc13799, \B_DOUT_TEMPR5[24] , 
        \B_DOUT_TEMPR5[23] , \B_DOUT_TEMPR5[22] , \B_DOUT_TEMPR5[21] , 
        \B_DOUT_TEMPR5[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2727 (.A(\B_DOUT_TEMPR111[12] ), .B(\B_DOUT_TEMPR112[12] ), 
        .C(\B_DOUT_TEMPR113[12] ), .D(\B_DOUT_TEMPR114[12] ), .Y(
        OR4_2727_Y));
    OR4 OR4_1621 (.A(\A_DOUT_TEMPR83[35] ), .B(\A_DOUT_TEMPR84[35] ), 
        .C(\A_DOUT_TEMPR85[35] ), .D(\A_DOUT_TEMPR86[35] ), .Y(
        OR4_1621_Y));
    OR4 OR4_636 (.A(OR4_1043_Y), .B(OR4_1832_Y), .C(OR4_913_Y), .D(
        OR4_1399_Y), .Y(OR4_636_Y));
    OR4 OR4_2521 (.A(\B_DOUT_TEMPR12[2] ), .B(\B_DOUT_TEMPR13[2] ), .C(
        \B_DOUT_TEMPR14[2] ), .D(\B_DOUT_TEMPR15[2] ), .Y(OR4_2521_Y));
    OR4 OR4_864 (.A(\A_DOUT_TEMPR32[19] ), .B(\A_DOUT_TEMPR33[19] ), 
        .C(\A_DOUT_TEMPR34[19] ), .D(\A_DOUT_TEMPR35[19] ), .Y(
        OR4_864_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%58%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R58C5 (
        .A_DOUT({nc13800, nc13801, nc13802, nc13803, nc13804, nc13805, 
        nc13806, nc13807, nc13808, nc13809, nc13810, nc13811, nc13812, 
        nc13813, nc13814, \A_DOUT_TEMPR58[29] , \A_DOUT_TEMPR58[28] , 
        \A_DOUT_TEMPR58[27] , \A_DOUT_TEMPR58[26] , 
        \A_DOUT_TEMPR58[25] }), .B_DOUT({nc13815, nc13816, nc13817, 
        nc13818, nc13819, nc13820, nc13821, nc13822, nc13823, nc13824, 
        nc13825, nc13826, nc13827, nc13828, nc13829, 
        \B_DOUT_TEMPR58[29] , \B_DOUT_TEMPR58[28] , 
        \B_DOUT_TEMPR58[27] , \B_DOUT_TEMPR58[26] , 
        \B_DOUT_TEMPR58[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[58][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1843 (.A(\A_DOUT_TEMPR48[29] ), .B(\A_DOUT_TEMPR49[29] ), 
        .C(\A_DOUT_TEMPR50[29] ), .D(\A_DOUT_TEMPR51[29] ), .Y(
        OR4_1843_Y));
    OR4 OR4_1723 (.A(\B_DOUT_TEMPR28[29] ), .B(\B_DOUT_TEMPR29[29] ), 
        .C(\B_DOUT_TEMPR30[29] ), .D(\B_DOUT_TEMPR31[29] ), .Y(
        OR4_1723_Y));
    OR4 OR4_562 (.A(\A_DOUT_TEMPR75[33] ), .B(\A_DOUT_TEMPR76[33] ), 
        .C(\A_DOUT_TEMPR77[33] ), .D(\A_DOUT_TEMPR78[33] ), .Y(
        OR4_562_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%100%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R100C0 (
        .A_DOUT({nc13830, nc13831, nc13832, nc13833, nc13834, nc13835, 
        nc13836, nc13837, nc13838, nc13839, nc13840, nc13841, nc13842, 
        nc13843, nc13844, \A_DOUT_TEMPR100[4] , \A_DOUT_TEMPR100[3] , 
        \A_DOUT_TEMPR100[2] , \A_DOUT_TEMPR100[1] , 
        \A_DOUT_TEMPR100[0] }), .B_DOUT({nc13845, nc13846, nc13847, 
        nc13848, nc13849, nc13850, nc13851, nc13852, nc13853, nc13854, 
        nc13855, nc13856, nc13857, nc13858, nc13859, 
        \B_DOUT_TEMPR100[4] , \B_DOUT_TEMPR100[3] , 
        \B_DOUT_TEMPR100[2] , \B_DOUT_TEMPR100[1] , 
        \B_DOUT_TEMPR100[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[100][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1125 (.A(\A_DOUT_TEMPR87[10] ), .B(\A_DOUT_TEMPR88[10] ), 
        .C(\A_DOUT_TEMPR89[10] ), .D(\A_DOUT_TEMPR90[10] ), .Y(
        OR4_1125_Y));
    OR4 OR4_742 (.A(\B_DOUT_TEMPR52[26] ), .B(\B_DOUT_TEMPR53[26] ), 
        .C(\B_DOUT_TEMPR54[26] ), .D(\B_DOUT_TEMPR55[26] ), .Y(
        OR4_742_Y));
    OR4 OR4_1550 (.A(\A_DOUT_TEMPR4[0] ), .B(\A_DOUT_TEMPR5[0] ), .C(
        \A_DOUT_TEMPR6[0] ), .D(\A_DOUT_TEMPR7[0] ), .Y(OR4_1550_Y));
    OR4 OR4_1394 (.A(\B_DOUT_TEMPR115[1] ), .B(\B_DOUT_TEMPR116[1] ), 
        .C(\B_DOUT_TEMPR117[1] ), .D(\B_DOUT_TEMPR118[1] ), .Y(
        OR4_1394_Y));
    OR4 OR4_1172 (.A(\A_DOUT_TEMPR32[28] ), .B(\A_DOUT_TEMPR33[28] ), 
        .C(\A_DOUT_TEMPR34[28] ), .D(\A_DOUT_TEMPR35[28] ), .Y(
        OR4_1172_Y));
    OR4 OR4_1749 (.A(\B_DOUT_TEMPR115[2] ), .B(\B_DOUT_TEMPR116[2] ), 
        .C(\B_DOUT_TEMPR117[2] ), .D(\B_DOUT_TEMPR118[2] ), .Y(
        OR4_1749_Y));
    OR4 OR4_346 (.A(\B_DOUT_TEMPR87[18] ), .B(\B_DOUT_TEMPR88[18] ), 
        .C(\B_DOUT_TEMPR89[18] ), .D(\B_DOUT_TEMPR90[18] ), .Y(
        OR4_346_Y));
    OR4 OR4_2318 (.A(OR4_804_Y), .B(OR4_1706_Y), .C(OR4_1379_Y), .D(
        OR4_2886_Y), .Y(OR4_2318_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%4%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R4C4 (
        .A_DOUT({nc13860, nc13861, nc13862, nc13863, nc13864, nc13865, 
        nc13866, nc13867, nc13868, nc13869, nc13870, nc13871, nc13872, 
        nc13873, nc13874, \A_DOUT_TEMPR4[24] , \A_DOUT_TEMPR4[23] , 
        \A_DOUT_TEMPR4[22] , \A_DOUT_TEMPR4[21] , \A_DOUT_TEMPR4[20] })
        , .B_DOUT({nc13875, nc13876, nc13877, nc13878, nc13879, 
        nc13880, nc13881, nc13882, nc13883, nc13884, nc13885, nc13886, 
        nc13887, nc13888, nc13889, \B_DOUT_TEMPR4[24] , 
        \B_DOUT_TEMPR4[23] , \B_DOUT_TEMPR4[22] , \B_DOUT_TEMPR4[21] , 
        \B_DOUT_TEMPR4[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1514 (.A(OR4_1001_Y), .B(OR4_775_Y), .C(OR4_1636_Y), .D(
        OR4_2866_Y), .Y(OR4_1514_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%106%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R106C6 (
        .A_DOUT({nc13890, nc13891, nc13892, nc13893, nc13894, nc13895, 
        nc13896, nc13897, nc13898, nc13899, nc13900, nc13901, nc13902, 
        nc13903, nc13904, \A_DOUT_TEMPR106[34] , \A_DOUT_TEMPR106[33] , 
        \A_DOUT_TEMPR106[32] , \A_DOUT_TEMPR106[31] , 
        \A_DOUT_TEMPR106[30] }), .B_DOUT({nc13905, nc13906, nc13907, 
        nc13908, nc13909, nc13910, nc13911, nc13912, nc13913, nc13914, 
        nc13915, nc13916, nc13917, nc13918, nc13919, 
        \B_DOUT_TEMPR106[34] , \B_DOUT_TEMPR106[33] , 
        \B_DOUT_TEMPR106[32] , \B_DOUT_TEMPR106[31] , 
        \B_DOUT_TEMPR106[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[106][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%51%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R51C7 (
        .A_DOUT({nc13920, nc13921, nc13922, nc13923, nc13924, nc13925, 
        nc13926, nc13927, nc13928, nc13929, nc13930, nc13931, nc13932, 
        nc13933, nc13934, \A_DOUT_TEMPR51[39] , \A_DOUT_TEMPR51[38] , 
        \A_DOUT_TEMPR51[37] , \A_DOUT_TEMPR51[36] , 
        \A_DOUT_TEMPR51[35] }), .B_DOUT({nc13935, nc13936, nc13937, 
        nc13938, nc13939, nc13940, nc13941, nc13942, nc13943, nc13944, 
        nc13945, nc13946, nc13947, nc13948, nc13949, 
        \B_DOUT_TEMPR51[39] , \B_DOUT_TEMPR51[38] , 
        \B_DOUT_TEMPR51[37] , \B_DOUT_TEMPR51[36] , 
        \B_DOUT_TEMPR51[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[51][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_547 (.A(\A_DOUT_TEMPR83[34] ), .B(\A_DOUT_TEMPR84[34] ), 
        .C(\A_DOUT_TEMPR85[34] ), .D(\A_DOUT_TEMPR86[34] ), .Y(
        OR4_547_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%75%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R75C2 (
        .A_DOUT({nc13950, nc13951, nc13952, nc13953, nc13954, nc13955, 
        nc13956, nc13957, nc13958, nc13959, nc13960, nc13961, nc13962, 
        nc13963, nc13964, \A_DOUT_TEMPR75[14] , \A_DOUT_TEMPR75[13] , 
        \A_DOUT_TEMPR75[12] , \A_DOUT_TEMPR75[11] , 
        \A_DOUT_TEMPR75[10] }), .B_DOUT({nc13965, nc13966, nc13967, 
        nc13968, nc13969, nc13970, nc13971, nc13972, nc13973, nc13974, 
        nc13975, nc13976, nc13977, nc13978, nc13979, 
        \B_DOUT_TEMPR75[14] , \B_DOUT_TEMPR75[13] , 
        \B_DOUT_TEMPR75[12] , \B_DOUT_TEMPR75[11] , 
        \B_DOUT_TEMPR75[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[75][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%87%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R87C5 (
        .A_DOUT({nc13980, nc13981, nc13982, nc13983, nc13984, nc13985, 
        nc13986, nc13987, nc13988, nc13989, nc13990, nc13991, nc13992, 
        nc13993, nc13994, \A_DOUT_TEMPR87[29] , \A_DOUT_TEMPR87[28] , 
        \A_DOUT_TEMPR87[27] , \A_DOUT_TEMPR87[26] , 
        \A_DOUT_TEMPR87[25] }), .B_DOUT({nc13995, nc13996, nc13997, 
        nc13998, nc13999, nc14000, nc14001, nc14002, nc14003, nc14004, 
        nc14005, nc14006, nc14007, nc14008, nc14009, 
        \B_DOUT_TEMPR87[29] , \B_DOUT_TEMPR87[28] , 
        \B_DOUT_TEMPR87[27] , \B_DOUT_TEMPR87[26] , 
        \B_DOUT_TEMPR87[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[87][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1146 (.A(\B_DOUT_TEMPR99[22] ), .B(\B_DOUT_TEMPR100[22] ), 
        .C(\B_DOUT_TEMPR101[22] ), .D(\B_DOUT_TEMPR102[22] ), .Y(
        OR4_1146_Y));
    OR4 OR4_1021 (.A(\B_DOUT_TEMPR79[8] ), .B(\B_DOUT_TEMPR80[8] ), .C(
        \B_DOUT_TEMPR81[8] ), .D(\B_DOUT_TEMPR82[8] ), .Y(OR4_1021_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%112%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R112C7 (
        .A_DOUT({nc14010, nc14011, nc14012, nc14013, nc14014, nc14015, 
        nc14016, nc14017, nc14018, nc14019, nc14020, nc14021, nc14022, 
        nc14023, nc14024, \A_DOUT_TEMPR112[39] , \A_DOUT_TEMPR112[38] , 
        \A_DOUT_TEMPR112[37] , \A_DOUT_TEMPR112[36] , 
        \A_DOUT_TEMPR112[35] }), .B_DOUT({nc14025, nc14026, nc14027, 
        nc14028, nc14029, nc14030, nc14031, nc14032, nc14033, nc14034, 
        nc14035, nc14036, nc14037, nc14038, nc14039, 
        \B_DOUT_TEMPR112[39] , \B_DOUT_TEMPR112[38] , 
        \B_DOUT_TEMPR112[37] , \B_DOUT_TEMPR112[36] , 
        \B_DOUT_TEMPR112[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[112][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2975 (.A(OR4_2869_Y), .B(OR4_798_Y), .C(OR4_1477_Y), .D(
        OR4_106_Y), .Y(OR4_2975_Y));
    OR4 OR4_1548 (.A(\A_DOUT_TEMPR12[3] ), .B(\A_DOUT_TEMPR13[3] ), .C(
        \A_DOUT_TEMPR14[3] ), .D(\A_DOUT_TEMPR15[3] ), .Y(OR4_1548_Y));
    OR4 OR4_134 (.A(\A_DOUT_TEMPR99[17] ), .B(\A_DOUT_TEMPR100[17] ), 
        .C(\A_DOUT_TEMPR101[17] ), .D(\A_DOUT_TEMPR102[17] ), .Y(
        OR4_134_Y));
    OR4 OR4_334 (.A(\B_DOUT_TEMPR44[1] ), .B(\B_DOUT_TEMPR45[1] ), .C(
        \B_DOUT_TEMPR46[1] ), .D(\B_DOUT_TEMPR47[1] ), .Y(OR4_334_Y));
    OR4 OR4_2299 (.A(OR4_2791_Y), .B(OR4_1916_Y), .C(OR4_354_Y), .D(
        OR4_1921_Y), .Y(OR4_2299_Y));
    OR4 OR4_457 (.A(\B_DOUT_TEMPR99[33] ), .B(\B_DOUT_TEMPR100[33] ), 
        .C(\B_DOUT_TEMPR101[33] ), .D(\B_DOUT_TEMPR102[33] ), .Y(
        OR4_457_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%7%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R7C1 (
        .A_DOUT({nc14040, nc14041, nc14042, nc14043, nc14044, nc14045, 
        nc14046, nc14047, nc14048, nc14049, nc14050, nc14051, nc14052, 
        nc14053, nc14054, \A_DOUT_TEMPR7[9] , \A_DOUT_TEMPR7[8] , 
        \A_DOUT_TEMPR7[7] , \A_DOUT_TEMPR7[6] , \A_DOUT_TEMPR7[5] }), 
        .B_DOUT({nc14055, nc14056, nc14057, nc14058, nc14059, nc14060, 
        nc14061, nc14062, nc14063, nc14064, nc14065, nc14066, nc14067, 
        nc14068, nc14069, \B_DOUT_TEMPR7[9] , \B_DOUT_TEMPR7[8] , 
        \B_DOUT_TEMPR7[7] , \B_DOUT_TEMPR7[6] , \B_DOUT_TEMPR7[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[7][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[1] , A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[1] , B_ADDR[13], B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2679 (.A(\B_DOUT_TEMPR12[20] ), .B(\B_DOUT_TEMPR13[20] ), 
        .C(\B_DOUT_TEMPR14[20] ), .D(\B_DOUT_TEMPR15[20] ), .Y(
        OR4_2679_Y));
    OR4 OR4_726 (.A(\B_DOUT_TEMPR44[7] ), .B(\B_DOUT_TEMPR45[7] ), .C(
        \B_DOUT_TEMPR46[7] ), .D(\B_DOUT_TEMPR47[7] ), .Y(OR4_726_Y));
    OR4 OR4_2554 (.A(\B_DOUT_TEMPR28[8] ), .B(\B_DOUT_TEMPR29[8] ), .C(
        \B_DOUT_TEMPR30[8] ), .D(\B_DOUT_TEMPR31[8] ), .Y(OR4_2554_Y));
    OR4 OR4_1211 (.A(\B_DOUT_TEMPR83[0] ), .B(\B_DOUT_TEMPR84[0] ), .C(
        \B_DOUT_TEMPR85[0] ), .D(\B_DOUT_TEMPR86[0] ), .Y(OR4_1211_Y));
    OR4 OR4_1955 (.A(\A_DOUT_TEMPR75[25] ), .B(\A_DOUT_TEMPR76[25] ), 
        .C(\A_DOUT_TEMPR77[25] ), .D(\A_DOUT_TEMPR78[25] ), .Y(
        OR4_1955_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%38%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R38C5 (
        .A_DOUT({nc14070, nc14071, nc14072, nc14073, nc14074, nc14075, 
        nc14076, nc14077, nc14078, nc14079, nc14080, nc14081, nc14082, 
        nc14083, nc14084, \A_DOUT_TEMPR38[29] , \A_DOUT_TEMPR38[28] , 
        \A_DOUT_TEMPR38[27] , \A_DOUT_TEMPR38[26] , 
        \A_DOUT_TEMPR38[25] }), .B_DOUT({nc14085, nc14086, nc14087, 
        nc14088, nc14089, nc14090, nc14091, nc14092, nc14093, nc14094, 
        nc14095, nc14096, nc14097, nc14098, nc14099, 
        \B_DOUT_TEMPR38[29] , \B_DOUT_TEMPR38[28] , 
        \B_DOUT_TEMPR38[27] , \B_DOUT_TEMPR38[26] , 
        \B_DOUT_TEMPR38[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[38][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1888 (.A(\A_DOUT_TEMPR12[16] ), .B(\A_DOUT_TEMPR13[16] ), 
        .C(\A_DOUT_TEMPR14[16] ), .D(\A_DOUT_TEMPR15[16] ), .Y(
        OR4_1888_Y));
    OR4 OR4_2289 (.A(\A_DOUT_TEMPR24[38] ), .B(\A_DOUT_TEMPR25[38] ), 
        .C(\A_DOUT_TEMPR26[38] ), .D(\A_DOUT_TEMPR27[38] ), .Y(
        OR4_2289_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%99%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R99C6 (
        .A_DOUT({nc14100, nc14101, nc14102, nc14103, nc14104, nc14105, 
        nc14106, nc14107, nc14108, nc14109, nc14110, nc14111, nc14112, 
        nc14113, nc14114, \A_DOUT_TEMPR99[34] , \A_DOUT_TEMPR99[33] , 
        \A_DOUT_TEMPR99[32] , \A_DOUT_TEMPR99[31] , 
        \A_DOUT_TEMPR99[30] }), .B_DOUT({nc14115, nc14116, nc14117, 
        nc14118, nc14119, nc14120, nc14121, nc14122, nc14123, nc14124, 
        nc14125, nc14126, nc14127, nc14128, nc14129, 
        \B_DOUT_TEMPR99[34] , \B_DOUT_TEMPR99[33] , 
        \B_DOUT_TEMPR99[32] , \B_DOUT_TEMPR99[31] , 
        \B_DOUT_TEMPR99[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[99][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2415 (.A(\A_DOUT_TEMPR48[18] ), .B(\A_DOUT_TEMPR49[18] ), 
        .C(\A_DOUT_TEMPR50[18] ), .D(\A_DOUT_TEMPR51[18] ), .Y(
        OR4_2415_Y));
    OR4 OR4_1659 (.A(\B_DOUT_TEMPR40[0] ), .B(\B_DOUT_TEMPR41[0] ), .C(
        \B_DOUT_TEMPR42[0] ), .D(\B_DOUT_TEMPR43[0] ), .Y(OR4_1659_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%29%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R29C3 (
        .A_DOUT({nc14130, nc14131, nc14132, nc14133, nc14134, nc14135, 
        nc14136, nc14137, nc14138, nc14139, nc14140, nc14141, nc14142, 
        nc14143, nc14144, \A_DOUT_TEMPR29[19] , \A_DOUT_TEMPR29[18] , 
        \A_DOUT_TEMPR29[17] , \A_DOUT_TEMPR29[16] , 
        \A_DOUT_TEMPR29[15] }), .B_DOUT({nc14145, nc14146, nc14147, 
        nc14148, nc14149, nc14150, nc14151, nc14152, nc14153, nc14154, 
        nc14155, nc14156, nc14157, nc14158, nc14159, 
        \B_DOUT_TEMPR29[19] , \B_DOUT_TEMPR29[18] , 
        \B_DOUT_TEMPR29[17] , \B_DOUT_TEMPR29[16] , 
        \B_DOUT_TEMPR29[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%85%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R85C7 (
        .A_DOUT({nc14160, nc14161, nc14162, nc14163, nc14164, nc14165, 
        nc14166, nc14167, nc14168, nc14169, nc14170, nc14171, nc14172, 
        nc14173, nc14174, \A_DOUT_TEMPR85[39] , \A_DOUT_TEMPR85[38] , 
        \A_DOUT_TEMPR85[37] , \A_DOUT_TEMPR85[36] , 
        \A_DOUT_TEMPR85[35] }), .B_DOUT({nc14175, nc14176, nc14177, 
        nc14178, nc14179, nc14180, nc14181, nc14182, nc14183, nc14184, 
        nc14185, nc14186, nc14187, nc14188, nc14189, 
        \B_DOUT_TEMPR85[39] , \B_DOUT_TEMPR85[38] , 
        \B_DOUT_TEMPR85[37] , \B_DOUT_TEMPR85[36] , 
        \B_DOUT_TEMPR85[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[85][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%66%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R66C1 (
        .A_DOUT({nc14190, nc14191, nc14192, nc14193, nc14194, nc14195, 
        nc14196, nc14197, nc14198, nc14199, nc14200, nc14201, nc14202, 
        nc14203, nc14204, \A_DOUT_TEMPR66[9] , \A_DOUT_TEMPR66[8] , 
        \A_DOUT_TEMPR66[7] , \A_DOUT_TEMPR66[6] , \A_DOUT_TEMPR66[5] })
        , .B_DOUT({nc14205, nc14206, nc14207, nc14208, nc14209, 
        nc14210, nc14211, nc14212, nc14213, nc14214, nc14215, nc14216, 
        nc14217, nc14218, nc14219, \B_DOUT_TEMPR66[9] , 
        \B_DOUT_TEMPR66[8] , \B_DOUT_TEMPR66[7] , \B_DOUT_TEMPR66[6] , 
        \B_DOUT_TEMPR66[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[66][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_521 (.A(OR4_3010_Y), .B(OR4_257_Y), .C(OR4_2955_Y), .D(
        OR4_273_Y), .Y(OR4_521_Y));
    OR4 OR4_528 (.A(\B_DOUT_TEMPR56[19] ), .B(\B_DOUT_TEMPR57[19] ), 
        .C(\B_DOUT_TEMPR58[19] ), .D(\B_DOUT_TEMPR59[19] ), .Y(
        OR4_528_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%31%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R31C7 (
        .A_DOUT({nc14220, nc14221, nc14222, nc14223, nc14224, nc14225, 
        nc14226, nc14227, nc14228, nc14229, nc14230, nc14231, nc14232, 
        nc14233, nc14234, \A_DOUT_TEMPR31[39] , \A_DOUT_TEMPR31[38] , 
        \A_DOUT_TEMPR31[37] , \A_DOUT_TEMPR31[36] , 
        \A_DOUT_TEMPR31[35] }), .B_DOUT({nc14235, nc14236, nc14237, 
        nc14238, nc14239, nc14240, nc14241, nc14242, nc14243, nc14244, 
        nc14245, nc14246, nc14247, nc14248, nc14249, 
        \B_DOUT_TEMPR31[39] , \B_DOUT_TEMPR31[38] , 
        \B_DOUT_TEMPR31[37] , \B_DOUT_TEMPR31[36] , 
        \B_DOUT_TEMPR31[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2251 (.A(\B_DOUT_TEMPR24[35] ), .B(\B_DOUT_TEMPR25[35] ), 
        .C(\B_DOUT_TEMPR26[35] ), .D(\B_DOUT_TEMPR27[35] ), .Y(
        OR4_2251_Y));
    OR4 OR4_1490 (.A(\B_DOUT_TEMPR83[5] ), .B(\B_DOUT_TEMPR84[5] ), .C(
        \B_DOUT_TEMPR85[5] ), .D(\B_DOUT_TEMPR86[5] ), .Y(OR4_1490_Y));
    OR4 OR4_2162 (.A(\A_DOUT_TEMPR60[26] ), .B(\A_DOUT_TEMPR61[26] ), 
        .C(\A_DOUT_TEMPR62[26] ), .D(\A_DOUT_TEMPR63[26] ), .Y(
        OR4_2162_Y));
    OR4 OR4_1009 (.A(\B_DOUT_TEMPR83[25] ), .B(\B_DOUT_TEMPR84[25] ), 
        .C(\B_DOUT_TEMPR85[25] ), .D(\B_DOUT_TEMPR86[25] ), .Y(
        OR4_1009_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%66%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R66C2 (
        .A_DOUT({nc14250, nc14251, nc14252, nc14253, nc14254, nc14255, 
        nc14256, nc14257, nc14258, nc14259, nc14260, nc14261, nc14262, 
        nc14263, nc14264, \A_DOUT_TEMPR66[14] , \A_DOUT_TEMPR66[13] , 
        \A_DOUT_TEMPR66[12] , \A_DOUT_TEMPR66[11] , 
        \A_DOUT_TEMPR66[10] }), .B_DOUT({nc14265, nc14266, nc14267, 
        nc14268, nc14269, nc14270, nc14271, nc14272, nc14273, nc14274, 
        nc14275, nc14276, nc14277, nc14278, nc14279, 
        \B_DOUT_TEMPR66[14] , \B_DOUT_TEMPR66[13] , 
        \B_DOUT_TEMPR66[12] , \B_DOUT_TEMPR66[11] , 
        \B_DOUT_TEMPR66[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[66][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2638 (.A(\A_DOUT_TEMPR99[29] ), .B(\A_DOUT_TEMPR100[29] ), 
        .C(\A_DOUT_TEMPR101[29] ), .D(\A_DOUT_TEMPR102[29] ), .Y(
        OR4_2638_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%27%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R27C3 (
        .A_DOUT({nc14280, nc14281, nc14282, nc14283, nc14284, nc14285, 
        nc14286, nc14287, nc14288, nc14289, nc14290, nc14291, nc14292, 
        nc14293, nc14294, \A_DOUT_TEMPR27[19] , \A_DOUT_TEMPR27[18] , 
        \A_DOUT_TEMPR27[17] , \A_DOUT_TEMPR27[16] , 
        \A_DOUT_TEMPR27[15] }), .B_DOUT({nc14295, nc14296, nc14297, 
        nc14298, nc14299, nc14300, nc14301, nc14302, nc14303, nc14304, 
        nc14305, nc14306, nc14307, nc14308, nc14309, 
        \B_DOUT_TEMPR27[19] , \B_DOUT_TEMPR27[18] , 
        \B_DOUT_TEMPR27[17] , \B_DOUT_TEMPR27[16] , 
        \B_DOUT_TEMPR27[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2716 (.A(OR4_849_Y), .B(OR4_1819_Y), .C(OR4_2507_Y), .D(
        OR4_1151_Y), .Y(OR4_2716_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%60%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R60C6 (
        .A_DOUT({nc14310, nc14311, nc14312, nc14313, nc14314, nc14315, 
        nc14316, nc14317, nc14318, nc14319, nc14320, nc14321, nc14322, 
        nc14323, nc14324, \A_DOUT_TEMPR60[34] , \A_DOUT_TEMPR60[33] , 
        \A_DOUT_TEMPR60[32] , \A_DOUT_TEMPR60[31] , 
        \A_DOUT_TEMPR60[30] }), .B_DOUT({nc14325, nc14326, nc14327, 
        nc14328, nc14329, nc14330, nc14331, nc14332, nc14333, nc14334, 
        nc14335, nc14336, nc14337, nc14338, nc14339, 
        \B_DOUT_TEMPR60[34] , \B_DOUT_TEMPR60[33] , 
        \B_DOUT_TEMPR60[32] , \B_DOUT_TEMPR60[31] , 
        \B_DOUT_TEMPR60[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[60][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%57%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R57C0 (
        .A_DOUT({nc14340, nc14341, nc14342, nc14343, nc14344, nc14345, 
        nc14346, nc14347, nc14348, nc14349, nc14350, nc14351, nc14352, 
        nc14353, nc14354, \A_DOUT_TEMPR57[4] , \A_DOUT_TEMPR57[3] , 
        \A_DOUT_TEMPR57[2] , \A_DOUT_TEMPR57[1] , \A_DOUT_TEMPR57[0] })
        , .B_DOUT({nc14355, nc14356, nc14357, nc14358, nc14359, 
        nc14360, nc14361, nc14362, nc14363, nc14364, nc14365, nc14366, 
        nc14367, nc14368, nc14369, \B_DOUT_TEMPR57[4] , 
        \B_DOUT_TEMPR57[3] , \B_DOUT_TEMPR57[2] , \B_DOUT_TEMPR57[1] , 
        \B_DOUT_TEMPR57[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[57][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1509 (.A(\A_DOUT_TEMPR68[11] ), .B(\A_DOUT_TEMPR69[11] ), 
        .C(\A_DOUT_TEMPR70[11] ), .D(\A_DOUT_TEMPR71[11] ), .Y(
        OR4_1509_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%60%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R60C5 (
        .A_DOUT({nc14370, nc14371, nc14372, nc14373, nc14374, nc14375, 
        nc14376, nc14377, nc14378, nc14379, nc14380, nc14381, nc14382, 
        nc14383, nc14384, \A_DOUT_TEMPR60[29] , \A_DOUT_TEMPR60[28] , 
        \A_DOUT_TEMPR60[27] , \A_DOUT_TEMPR60[26] , 
        \A_DOUT_TEMPR60[25] }), .B_DOUT({nc14385, nc14386, nc14387, 
        nc14388, nc14389, nc14390, nc14391, nc14392, nc14393, nc14394, 
        nc14395, nc14396, nc14397, nc14398, nc14399, 
        \B_DOUT_TEMPR60[29] , \B_DOUT_TEMPR60[28] , 
        \B_DOUT_TEMPR60[27] , \B_DOUT_TEMPR60[26] , 
        \B_DOUT_TEMPR60[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[60][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%118%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R118C4 (
        .A_DOUT({nc14400, nc14401, nc14402, nc14403, nc14404, nc14405, 
        nc14406, nc14407, nc14408, nc14409, nc14410, nc14411, nc14412, 
        nc14413, nc14414, \A_DOUT_TEMPR118[24] , \A_DOUT_TEMPR118[23] , 
        \A_DOUT_TEMPR118[22] , \A_DOUT_TEMPR118[21] , 
        \A_DOUT_TEMPR118[20] }), .B_DOUT({nc14415, nc14416, nc14417, 
        nc14418, nc14419, nc14420, nc14421, nc14422, nc14423, nc14424, 
        nc14425, nc14426, nc14427, nc14428, nc14429, 
        \B_DOUT_TEMPR118[24] , \B_DOUT_TEMPR118[23] , 
        \B_DOUT_TEMPR118[22] , \B_DOUT_TEMPR118[21] , 
        \B_DOUT_TEMPR118[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[118][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1638 (.A(\A_DOUT_TEMPR56[18] ), .B(\A_DOUT_TEMPR57[18] ), 
        .C(\A_DOUT_TEMPR58[18] ), .D(\A_DOUT_TEMPR59[18] ), .Y(
        OR4_1638_Y));
    OR4 OR4_836 (.A(\A_DOUT_TEMPR28[29] ), .B(\A_DOUT_TEMPR29[29] ), 
        .C(\A_DOUT_TEMPR30[29] ), .D(\A_DOUT_TEMPR31[29] ), .Y(
        OR4_836_Y));
    OR4 OR4_325 (.A(\B_DOUT_TEMPR44[8] ), .B(\B_DOUT_TEMPR45[8] ), .C(
        \B_DOUT_TEMPR46[8] ), .D(\B_DOUT_TEMPR47[8] ), .Y(OR4_325_Y));
    OR4 OR4_1279 (.A(OR4_629_Y), .B(OR4_2420_Y), .C(OR4_887_Y), .D(
        OR4_2421_Y), .Y(OR4_1279_Y));
    OR4 OR4_57 (.A(OR4_1970_Y), .B(OR4_117_Y), .C(OR4_1191_Y), .D(
        OR4_936_Y), .Y(OR4_57_Y));
    OR4 OR4_2828 (.A(\A_DOUT_TEMPR56[10] ), .B(\A_DOUT_TEMPR57[10] ), 
        .C(\A_DOUT_TEMPR58[10] ), .D(\A_DOUT_TEMPR59[10] ), .Y(
        OR4_2828_Y));
    OR4 OR4_746 (.A(\B_DOUT_TEMPR16[18] ), .B(\B_DOUT_TEMPR17[18] ), 
        .C(\B_DOUT_TEMPR18[18] ), .D(\B_DOUT_TEMPR19[18] ), .Y(
        OR4_746_Y));
    OR4 OR4_1295 (.A(OR4_3005_Y), .B(OR4_971_Y), .C(OR4_1619_Y), .D(
        OR4_243_Y), .Y(OR4_1295_Y));
    OR4 OR4_1544 (.A(\B_DOUT_TEMPR115[34] ), .B(\B_DOUT_TEMPR116[34] ), 
        .C(\B_DOUT_TEMPR117[34] ), .D(\B_DOUT_TEMPR118[34] ), .Y(
        OR4_1544_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%97%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R97C1 (
        .A_DOUT({nc14430, nc14431, nc14432, nc14433, nc14434, nc14435, 
        nc14436, nc14437, nc14438, nc14439, nc14440, nc14441, nc14442, 
        nc14443, nc14444, \A_DOUT_TEMPR97[9] , \A_DOUT_TEMPR97[8] , 
        \A_DOUT_TEMPR97[7] , \A_DOUT_TEMPR97[6] , \A_DOUT_TEMPR97[5] })
        , .B_DOUT({nc14445, nc14446, nc14447, nc14448, nc14449, 
        nc14450, nc14451, nc14452, nc14453, nc14454, nc14455, nc14456, 
        nc14457, nc14458, nc14459, \B_DOUT_TEMPR97[9] , 
        \B_DOUT_TEMPR97[8] , \B_DOUT_TEMPR97[7] , \B_DOUT_TEMPR97[6] , 
        \B_DOUT_TEMPR97[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[97][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1064 (.A(\A_DOUT_TEMPR44[17] ), .B(\A_DOUT_TEMPR45[17] ), 
        .C(\A_DOUT_TEMPR46[17] ), .D(\A_DOUT_TEMPR47[17] ), .Y(
        OR4_1064_Y));
    OR4 OR4_330 (.A(\A_DOUT_TEMPR95[17] ), .B(\A_DOUT_TEMPR96[17] ), 
        .C(\A_DOUT_TEMPR97[17] ), .D(\A_DOUT_TEMPR98[17] ), .Y(
        OR4_330_Y));
    OR4 OR4_2701 (.A(\B_DOUT_TEMPR44[31] ), .B(\B_DOUT_TEMPR45[31] ), 
        .C(\B_DOUT_TEMPR46[31] ), .D(\B_DOUT_TEMPR47[31] ), .Y(
        OR4_2701_Y));
    OR4 OR4_1066 (.A(\A_DOUT_TEMPR24[39] ), .B(\A_DOUT_TEMPR25[39] ), 
        .C(\A_DOUT_TEMPR26[39] ), .D(\A_DOUT_TEMPR27[39] ), .Y(
        OR4_1066_Y));
    OR4 OR4_1788 (.A(\B_DOUT_TEMPR107[30] ), .B(\B_DOUT_TEMPR108[30] ), 
        .C(\B_DOUT_TEMPR109[30] ), .D(\B_DOUT_TEMPR110[30] ), .Y(
        OR4_1788_Y));
    OR4 OR4_1302 (.A(\A_DOUT_TEMPR91[38] ), .B(\A_DOUT_TEMPR92[38] ), 
        .C(\A_DOUT_TEMPR93[38] ), .D(\A_DOUT_TEMPR94[38] ), .Y(
        OR4_1302_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%72%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R72C5 (
        .A_DOUT({nc14460, nc14461, nc14462, nc14463, nc14464, nc14465, 
        nc14466, nc14467, nc14468, nc14469, nc14470, nc14471, nc14472, 
        nc14473, nc14474, \A_DOUT_TEMPR72[29] , \A_DOUT_TEMPR72[28] , 
        \A_DOUT_TEMPR72[27] , \A_DOUT_TEMPR72[26] , 
        \A_DOUT_TEMPR72[25] }), .B_DOUT({nc14475, nc14476, nc14477, 
        nc14478, nc14479, nc14480, nc14481, nc14482, nc14483, nc14484, 
        nc14485, nc14486, nc14487, nc14488, nc14489, 
        \B_DOUT_TEMPR72[29] , \B_DOUT_TEMPR72[28] , 
        \B_DOUT_TEMPR72[27] , \B_DOUT_TEMPR72[26] , 
        \B_DOUT_TEMPR72[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[72][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2077 (.A(\B_DOUT_TEMPR75[26] ), .B(\B_DOUT_TEMPR76[26] ), 
        .C(\B_DOUT_TEMPR77[26] ), .D(\B_DOUT_TEMPR78[26] ), .Y(
        OR4_2077_Y));
    OR4 OR4_180 (.A(OR4_504_Y), .B(OR4_3027_Y), .C(OR4_1317_Y), .D(
        OR4_2210_Y), .Y(OR4_180_Y));
    OR4 OR4_2379 (.A(\B_DOUT_TEMPR68[19] ), .B(\B_DOUT_TEMPR69[19] ), 
        .C(\B_DOUT_TEMPR70[19] ), .D(\B_DOUT_TEMPR71[19] ), .Y(
        OR4_2379_Y));
    OR4 OR4_2277 (.A(OR4_2370_Y), .B(OR4_249_Y), .C(OR4_2965_Y), .D(
        OR4_1409_Y), .Y(OR4_2277_Y));
    OR4 OR4_497 (.A(OR4_1531_Y), .B(OR4_2338_Y), .C(OR2_33_Y), .D(
        \B_DOUT_TEMPR74[28] ), .Y(OR4_497_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[17]  (.A(CFG3_8_Y), .B(
        CFG3_21_Y), .Y(\BLKY2[17] ));
    OR4 OR4_1363 (.A(\B_DOUT_TEMPR28[9] ), .B(\B_DOUT_TEMPR29[9] ), .C(
        \B_DOUT_TEMPR30[9] ), .D(\B_DOUT_TEMPR31[9] ), .Y(OR4_1363_Y));
    OR4 OR4_2148 (.A(OR4_2515_Y), .B(OR4_918_Y), .C(OR2_13_Y), .D(
        \A_DOUT_TEMPR74[3] ), .Y(OR4_2148_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%72%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R72C1 (
        .A_DOUT({nc14490, nc14491, nc14492, nc14493, nc14494, nc14495, 
        nc14496, nc14497, nc14498, nc14499, nc14500, nc14501, nc14502, 
        nc14503, nc14504, \A_DOUT_TEMPR72[9] , \A_DOUT_TEMPR72[8] , 
        \A_DOUT_TEMPR72[7] , \A_DOUT_TEMPR72[6] , \A_DOUT_TEMPR72[5] })
        , .B_DOUT({nc14505, nc14506, nc14507, nc14508, nc14509, 
        nc14510, nc14511, nc14512, nc14513, nc14514, nc14515, nc14516, 
        nc14517, nc14518, nc14519, \B_DOUT_TEMPR72[9] , 
        \B_DOUT_TEMPR72[8] , \B_DOUT_TEMPR72[7] , \B_DOUT_TEMPR72[6] , 
        \B_DOUT_TEMPR72[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[72][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[19]  (.A(CFG3_20_Y), .B(
        CFG3_21_Y), .Y(\BLKY2[19] ));
    OR4 OR4_541 (.A(\A_DOUT_TEMPR64[34] ), .B(\A_DOUT_TEMPR65[34] ), 
        .C(\A_DOUT_TEMPR66[34] ), .D(\A_DOUT_TEMPR67[34] ), .Y(
        OR4_541_Y));
    OR4 OR4_548 (.A(\B_DOUT_TEMPR60[30] ), .B(\B_DOUT_TEMPR61[30] ), 
        .C(\B_DOUT_TEMPR62[30] ), .D(\B_DOUT_TEMPR63[30] ), .Y(
        OR4_548_Y));
    OR4 OR4_820 (.A(\B_DOUT_TEMPR4[4] ), .B(\B_DOUT_TEMPR5[4] ), .C(
        \B_DOUT_TEMPR6[4] ), .D(\B_DOUT_TEMPR7[4] ), .Y(OR4_820_Y));
    OR4 OR4_2970 (.A(OR4_1739_Y), .B(OR4_1563_Y), .C(OR4_1504_Y), .D(
        OR4_1223_Y), .Y(OR4_2970_Y));
    OR4 OR4_1241 (.A(\A_DOUT_TEMPR68[13] ), .B(\A_DOUT_TEMPR69[13] ), 
        .C(\A_DOUT_TEMPR70[13] ), .D(\A_DOUT_TEMPR71[13] ), .Y(
        OR4_1241_Y));
    OR4 OR4_688 (.A(\B_DOUT_TEMPR56[3] ), .B(\B_DOUT_TEMPR57[3] ), .C(
        \B_DOUT_TEMPR58[3] ), .D(\B_DOUT_TEMPR59[3] ), .Y(OR4_688_Y));
    OR4 OR4_520 (.A(\B_DOUT_TEMPR8[8] ), .B(\B_DOUT_TEMPR9[8] ), .C(
        \B_DOUT_TEMPR10[8] ), .D(\B_DOUT_TEMPR11[8] ), .Y(OR4_520_Y));
    OR4 OR4_1057 (.A(\B_DOUT_TEMPR28[15] ), .B(\B_DOUT_TEMPR29[15] ), 
        .C(\B_DOUT_TEMPR30[15] ), .D(\B_DOUT_TEMPR31[15] ), .Y(
        OR4_1057_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%87%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R87C2 (
        .A_DOUT({nc14520, nc14521, nc14522, nc14523, nc14524, nc14525, 
        nc14526, nc14527, nc14528, nc14529, nc14530, nc14531, nc14532, 
        nc14533, nc14534, \A_DOUT_TEMPR87[14] , \A_DOUT_TEMPR87[13] , 
        \A_DOUT_TEMPR87[12] , \A_DOUT_TEMPR87[11] , 
        \A_DOUT_TEMPR87[10] }), .B_DOUT({nc14535, nc14536, nc14537, 
        nc14538, nc14539, nc14540, nc14541, nc14542, nc14543, nc14544, 
        nc14545, nc14546, nc14547, nc14548, nc14549, 
        \B_DOUT_TEMPR87[14] , \B_DOUT_TEMPR87[13] , 
        \B_DOUT_TEMPR87[12] , \B_DOUT_TEMPR87[11] , 
        \B_DOUT_TEMPR87[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[87][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[13]  (.A(CFG3_1_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[13] ));
    OR4 OR4_1359 (.A(\B_DOUT_TEMPR16[10] ), .B(\B_DOUT_TEMPR17[10] ), 
        .C(\B_DOUT_TEMPR18[10] ), .D(\B_DOUT_TEMPR19[10] ), .Y(
        OR4_1359_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[15]  (.A(CFG3_2_Y), .B(
        CFG3_15_Y), .Y(\BLKY2[15] ));
    OR4 OR4_1505 (.A(\A_DOUT_TEMPR64[19] ), .B(\A_DOUT_TEMPR65[19] ), 
        .C(\A_DOUT_TEMPR66[19] ), .D(\A_DOUT_TEMPR67[19] ), .Y(
        OR4_1505_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[22]  (.A(CFG3_19_Y), .B(
        CFG3_21_Y), .Y(\BLKY2[22] ));
    OR4 OR4_1257 (.A(\B_DOUT_TEMPR103[27] ), .B(\B_DOUT_TEMPR104[27] ), 
        .C(\B_DOUT_TEMPR105[27] ), .D(\B_DOUT_TEMPR106[27] ), .Y(
        OR4_1257_Y));
    OR2 OR2_57 (.A(\B_DOUT_TEMPR72[32] ), .B(\B_DOUT_TEMPR73[32] ), .Y(
        OR2_57_Y));
    OR4 OR4_50 (.A(\B_DOUT_TEMPR52[17] ), .B(\B_DOUT_TEMPR53[17] ), .C(
        \B_DOUT_TEMPR54[17] ), .D(\B_DOUT_TEMPR55[17] ), .Y(OR4_50_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%101%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R101C0 (
        .A_DOUT({nc14550, nc14551, nc14552, nc14553, nc14554, nc14555, 
        nc14556, nc14557, nc14558, nc14559, nc14560, nc14561, nc14562, 
        nc14563, nc14564, \A_DOUT_TEMPR101[4] , \A_DOUT_TEMPR101[3] , 
        \A_DOUT_TEMPR101[2] , \A_DOUT_TEMPR101[1] , 
        \A_DOUT_TEMPR101[0] }), .B_DOUT({nc14565, nc14566, nc14567, 
        nc14568, nc14569, nc14570, nc14571, nc14572, nc14573, nc14574, 
        nc14575, nc14576, nc14577, nc14578, nc14579, 
        \B_DOUT_TEMPR101[4] , \B_DOUT_TEMPR101[3] , 
        \B_DOUT_TEMPR101[2] , \B_DOUT_TEMPR101[1] , 
        \B_DOUT_TEMPR101[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[101][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2843 (.A(\B_DOUT_TEMPR40[25] ), .B(\B_DOUT_TEMPR41[25] ), 
        .C(\B_DOUT_TEMPR42[25] ), .D(\B_DOUT_TEMPR43[25] ), .Y(
        OR4_2843_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%37%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R37C0 (
        .A_DOUT({nc14580, nc14581, nc14582, nc14583, nc14584, nc14585, 
        nc14586, nc14587, nc14588, nc14589, nc14590, nc14591, nc14592, 
        nc14593, nc14594, \A_DOUT_TEMPR37[4] , \A_DOUT_TEMPR37[3] , 
        \A_DOUT_TEMPR37[2] , \A_DOUT_TEMPR37[1] , \A_DOUT_TEMPR37[0] })
        , .B_DOUT({nc14595, nc14596, nc14597, nc14598, nc14599, 
        nc14600, nc14601, nc14602, nc14603, nc14604, nc14605, nc14606, 
        nc14607, nc14608, nc14609, \B_DOUT_TEMPR37[4] , 
        \B_DOUT_TEMPR37[3] , \B_DOUT_TEMPR37[2] , \B_DOUT_TEMPR37[1] , 
        \B_DOUT_TEMPR37[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[37][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%43%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R43C5 (
        .A_DOUT({nc14610, nc14611, nc14612, nc14613, nc14614, nc14615, 
        nc14616, nc14617, nc14618, nc14619, nc14620, nc14621, nc14622, 
        nc14623, nc14624, \A_DOUT_TEMPR43[29] , \A_DOUT_TEMPR43[28] , 
        \A_DOUT_TEMPR43[27] , \A_DOUT_TEMPR43[26] , 
        \A_DOUT_TEMPR43[25] }), .B_DOUT({nc14625, nc14626, nc14627, 
        nc14628, nc14629, nc14630, nc14631, nc14632, nc14633, nc14634, 
        nc14635, nc14636, nc14637, nc14638, nc14639, 
        \B_DOUT_TEMPR43[29] , \B_DOUT_TEMPR43[28] , 
        \B_DOUT_TEMPR43[27] , \B_DOUT_TEMPR43[26] , 
        \B_DOUT_TEMPR43[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[43][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2403 (.A(\B_DOUT_TEMPR91[18] ), .B(\B_DOUT_TEMPR92[18] ), 
        .C(\B_DOUT_TEMPR93[18] ), .D(\B_DOUT_TEMPR94[18] ), .Y(
        OR4_2403_Y));
    OR4 OR4_2728 (.A(\A_DOUT_TEMPR24[35] ), .B(\A_DOUT_TEMPR25[35] ), 
        .C(\A_DOUT_TEMPR26[35] ), .D(\A_DOUT_TEMPR27[35] ), .Y(
        OR4_2728_Y));
    OR4 OR4_724 (.A(\B_DOUT_TEMPR111[0] ), .B(\B_DOUT_TEMPR112[0] ), 
        .C(\B_DOUT_TEMPR113[0] ), .D(\B_DOUT_TEMPR114[0] ), .Y(
        OR4_724_Y));
    OR4 OR4_1950 (.A(\A_DOUT_TEMPR75[0] ), .B(\A_DOUT_TEMPR76[0] ), .C(
        \A_DOUT_TEMPR77[0] ), .D(\A_DOUT_TEMPR78[0] ), .Y(OR4_1950_Y));
    OR4 OR4_981 (.A(\B_DOUT_TEMPR91[38] ), .B(\B_DOUT_TEMPR92[38] ), 
        .C(\B_DOUT_TEMPR93[38] ), .D(\B_DOUT_TEMPR94[38] ), .Y(
        OR4_981_Y));
    OR4 OR4_345 (.A(OR4_1455_Y), .B(OR4_2664_Y), .C(OR2_20_Y), .D(
        \B_DOUT_TEMPR74[11] ), .Y(OR4_345_Y));
    OR4 OR4_2749 (.A(\A_DOUT_TEMPR107[1] ), .B(\A_DOUT_TEMPR108[1] ), 
        .C(\A_DOUT_TEMPR109[1] ), .D(\A_DOUT_TEMPR110[1] ), .Y(
        OR4_2749_Y));
    OR4 \OR4_A_DOUT[20]  (.A(OR4_178_Y), .B(OR4_2471_Y), .C(OR4_2671_Y)
        , .D(OR4_1013_Y), .Y(A_DOUT[20]));
    OR4 OR4_2772 (.A(\A_DOUT_TEMPR64[31] ), .B(\A_DOUT_TEMPR65[31] ), 
        .C(\A_DOUT_TEMPR66[31] ), .D(\A_DOUT_TEMPR67[31] ), .Y(
        OR4_2772_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%68%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R68C5 (
        .A_DOUT({nc14640, nc14641, nc14642, nc14643, nc14644, nc14645, 
        nc14646, nc14647, nc14648, nc14649, nc14650, nc14651, nc14652, 
        nc14653, nc14654, \A_DOUT_TEMPR68[29] , \A_DOUT_TEMPR68[28] , 
        \A_DOUT_TEMPR68[27] , \A_DOUT_TEMPR68[26] , 
        \A_DOUT_TEMPR68[25] }), .B_DOUT({nc14655, nc14656, nc14657, 
        nc14658, nc14659, nc14660, nc14661, nc14662, nc14663, nc14664, 
        nc14665, nc14666, nc14667, nc14668, nc14669, 
        \B_DOUT_TEMPR68[29] , \B_DOUT_TEMPR68[28] , 
        \B_DOUT_TEMPR68[27] , \B_DOUT_TEMPR68[26] , 
        \B_DOUT_TEMPR68[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[68][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%111%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R111C4 (
        .A_DOUT({nc14670, nc14671, nc14672, nc14673, nc14674, nc14675, 
        nc14676, nc14677, nc14678, nc14679, nc14680, nc14681, nc14682, 
        nc14683, nc14684, \A_DOUT_TEMPR111[24] , \A_DOUT_TEMPR111[23] , 
        \A_DOUT_TEMPR111[22] , \A_DOUT_TEMPR111[21] , 
        \A_DOUT_TEMPR111[20] }), .B_DOUT({nc14685, nc14686, nc14687, 
        nc14688, nc14689, nc14690, nc14691, nc14692, nc14693, nc14694, 
        nc14695, nc14696, nc14697, nc14698, nc14699, 
        \B_DOUT_TEMPR111[24] , \B_DOUT_TEMPR111[23] , 
        \B_DOUT_TEMPR111[22] , \B_DOUT_TEMPR111[21] , 
        \B_DOUT_TEMPR111[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[111][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%29%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R29C5 (
        .A_DOUT({nc14700, nc14701, nc14702, nc14703, nc14704, nc14705, 
        nc14706, nc14707, nc14708, nc14709, nc14710, nc14711, nc14712, 
        nc14713, nc14714, \A_DOUT_TEMPR29[29] , \A_DOUT_TEMPR29[28] , 
        \A_DOUT_TEMPR29[27] , \A_DOUT_TEMPR29[26] , 
        \A_DOUT_TEMPR29[25] }), .B_DOUT({nc14715, nc14716, nc14717, 
        nc14718, nc14719, nc14720, nc14721, nc14722, nc14723, nc14724, 
        nc14725, nc14726, nc14727, nc14728, nc14729, 
        \B_DOUT_TEMPR29[29] , \B_DOUT_TEMPR29[28] , 
        \B_DOUT_TEMPR29[27] , \B_DOUT_TEMPR29[26] , 
        \B_DOUT_TEMPR29[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%26%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R26C5 (
        .A_DOUT({nc14730, nc14731, nc14732, nc14733, nc14734, nc14735, 
        nc14736, nc14737, nc14738, nc14739, nc14740, nc14741, nc14742, 
        nc14743, nc14744, \A_DOUT_TEMPR26[29] , \A_DOUT_TEMPR26[28] , 
        \A_DOUT_TEMPR26[27] , \A_DOUT_TEMPR26[26] , 
        \A_DOUT_TEMPR26[25] }), .B_DOUT({nc14745, nc14746, nc14747, 
        nc14748, nc14749, nc14750, nc14751, nc14752, nc14753, nc14754, 
        nc14755, nc14756, nc14757, nc14758, nc14759, 
        \B_DOUT_TEMPR26[29] , \B_DOUT_TEMPR26[28] , 
        \B_DOUT_TEMPR26[27] , \B_DOUT_TEMPR26[26] , 
        \B_DOUT_TEMPR26[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%3%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R3C1 (
        .A_DOUT({nc14760, nc14761, nc14762, nc14763, nc14764, nc14765, 
        nc14766, nc14767, nc14768, nc14769, nc14770, nc14771, nc14772, 
        nc14773, nc14774, \A_DOUT_TEMPR3[9] , \A_DOUT_TEMPR3[8] , 
        \A_DOUT_TEMPR3[7] , \A_DOUT_TEMPR3[6] , \A_DOUT_TEMPR3[5] }), 
        .B_DOUT({nc14775, nc14776, nc14777, nc14778, nc14779, nc14780, 
        nc14781, nc14782, nc14783, nc14784, nc14785, nc14786, nc14787, 
        nc14788, nc14789, \B_DOUT_TEMPR3[9] , \B_DOUT_TEMPR3[8] , 
        \B_DOUT_TEMPR3[7] , \B_DOUT_TEMPR3[6] , \B_DOUT_TEMPR3[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[3][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[0] , A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[0] , B_ADDR[13], B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%0%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R0C1 (
        .A_DOUT({nc14790, nc14791, nc14792, nc14793, nc14794, nc14795, 
        nc14796, nc14797, nc14798, nc14799, nc14800, nc14801, nc14802, 
        nc14803, nc14804, \A_DOUT_TEMPR0[9] , \A_DOUT_TEMPR0[8] , 
        \A_DOUT_TEMPR0[7] , \A_DOUT_TEMPR0[6] , \A_DOUT_TEMPR0[5] }), 
        .B_DOUT({nc14805, nc14806, nc14807, nc14808, nc14809, nc14810, 
        nc14811, nc14812, nc14813, nc14814, nc14815, nc14816, nc14817, 
        nc14818, nc14819, \B_DOUT_TEMPR0[9] , \B_DOUT_TEMPR0[8] , 
        \B_DOUT_TEMPR0[7] , \B_DOUT_TEMPR0[6] , \B_DOUT_TEMPR0[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[0][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_672 (.A(\A_DOUT_TEMPR52[23] ), .B(\A_DOUT_TEMPR53[23] ), 
        .C(\A_DOUT_TEMPR54[23] ), .D(\A_DOUT_TEMPR55[23] ), .Y(
        OR4_672_Y));
    OR4 OR4_2517 (.A(\A_DOUT_TEMPR115[24] ), .B(\A_DOUT_TEMPR116[24] ), 
        .C(\A_DOUT_TEMPR117[24] ), .D(\A_DOUT_TEMPR118[24] ), .Y(
        OR4_2517_Y));
    OR4 OR4_418 (.A(\A_DOUT_TEMPR103[6] ), .B(\A_DOUT_TEMPR104[6] ), 
        .C(\A_DOUT_TEMPR105[6] ), .D(\A_DOUT_TEMPR106[6] ), .Y(
        OR4_418_Y));
    OR4 OR4_2269 (.A(\B_DOUT_TEMPR52[18] ), .B(\B_DOUT_TEMPR53[18] ), 
        .C(\B_DOUT_TEMPR54[18] ), .D(\B_DOUT_TEMPR55[18] ), .Y(
        OR4_2269_Y));
    OR4 OR4_1696 (.A(OR4_2139_Y), .B(OR4_36_Y), .C(OR4_2738_Y), .D(
        OR4_1193_Y), .Y(OR4_1696_Y));
    OR4 OR4_2146 (.A(\A_DOUT_TEMPR0[3] ), .B(\A_DOUT_TEMPR1[3] ), .C(
        \A_DOUT_TEMPR2[3] ), .D(\A_DOUT_TEMPR3[3] ), .Y(OR4_2146_Y));
    OR4 OR4_2991 (.A(OR4_712_Y), .B(OR4_1624_Y), .C(OR4_1292_Y), .D(
        OR4_2803_Y), .Y(OR4_2991_Y));
    OR4 OR4_514 (.A(\A_DOUT_TEMPR44[38] ), .B(\A_DOUT_TEMPR45[38] ), 
        .C(\A_DOUT_TEMPR46[38] ), .D(\A_DOUT_TEMPR47[38] ), .Y(
        OR4_514_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%16%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R16C1 (
        .A_DOUT({nc14820, nc14821, nc14822, nc14823, nc14824, nc14825, 
        nc14826, nc14827, nc14828, nc14829, nc14830, nc14831, nc14832, 
        nc14833, nc14834, \A_DOUT_TEMPR16[9] , \A_DOUT_TEMPR16[8] , 
        \A_DOUT_TEMPR16[7] , \A_DOUT_TEMPR16[6] , \A_DOUT_TEMPR16[5] })
        , .B_DOUT({nc14835, nc14836, nc14837, nc14838, nc14839, 
        nc14840, nc14841, nc14842, nc14843, nc14844, nc14845, nc14846, 
        nc14847, nc14848, nc14849, \B_DOUT_TEMPR16[9] , 
        \B_DOUT_TEMPR16[8] , \B_DOUT_TEMPR16[7] , \B_DOUT_TEMPR16[6] , 
        \B_DOUT_TEMPR16[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1190 (.A(\A_DOUT_TEMPR64[37] ), .B(\A_DOUT_TEMPR65[37] ), 
        .C(\A_DOUT_TEMPR66[37] ), .D(\A_DOUT_TEMPR67[37] ), .Y(
        OR4_1190_Y));
    OR4 OR4_2548 (.A(\A_DOUT_TEMPR107[23] ), .B(\A_DOUT_TEMPR108[23] ), 
        .C(\A_DOUT_TEMPR109[23] ), .D(\A_DOUT_TEMPR110[23] ), .Y(
        OR4_2548_Y));
    OR4 OR4_927 (.A(OR4_677_Y), .B(OR4_2095_Y), .C(OR4_1586_Y), .D(
        OR4_1569_Y), .Y(OR4_927_Y));
    OR4 OR4_234 (.A(\B_DOUT_TEMPR48[33] ), .B(\B_DOUT_TEMPR49[33] ), 
        .C(\B_DOUT_TEMPR50[33] ), .D(\B_DOUT_TEMPR51[33] ), .Y(
        OR4_234_Y));
    OR4 OR4_2839 (.A(\A_DOUT_TEMPR20[11] ), .B(\A_DOUT_TEMPR21[11] ), 
        .C(\A_DOUT_TEMPR22[11] ), .D(\A_DOUT_TEMPR23[11] ), .Y(
        OR4_2839_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%46%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R46C4 (
        .A_DOUT({nc14850, nc14851, nc14852, nc14853, nc14854, nc14855, 
        nc14856, nc14857, nc14858, nc14859, nc14860, nc14861, nc14862, 
        nc14863, nc14864, \A_DOUT_TEMPR46[24] , \A_DOUT_TEMPR46[23] , 
        \A_DOUT_TEMPR46[22] , \A_DOUT_TEMPR46[21] , 
        \A_DOUT_TEMPR46[20] }), .B_DOUT({nc14865, nc14866, nc14867, 
        nc14868, nc14869, nc14870, nc14871, nc14872, nc14873, nc14874, 
        nc14875, nc14876, nc14877, nc14878, nc14879, 
        \B_DOUT_TEMPR46[24] , \B_DOUT_TEMPR46[23] , 
        \B_DOUT_TEMPR46[22] , \B_DOUT_TEMPR46[21] , 
        \B_DOUT_TEMPR46[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[46][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[16]  (.A(CFG3_17_Y), .B(
        CFG3_3_Y), .Y(\BLKX2[16] ));
    OR4 OR4_1908 (.A(OR4_1199_Y), .B(OR4_2358_Y), .C(OR2_12_Y), .D(
        \B_DOUT_TEMPR74[14] ), .Y(OR4_1908_Y));
    OR4 OR4_1752 (.A(\B_DOUT_TEMPR28[39] ), .B(\B_DOUT_TEMPR29[39] ), 
        .C(\B_DOUT_TEMPR30[39] ), .D(\B_DOUT_TEMPR31[39] ), .Y(
        OR4_1752_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%61%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R61C7 (
        .A_DOUT({nc14880, nc14881, nc14882, nc14883, nc14884, nc14885, 
        nc14886, nc14887, nc14888, nc14889, nc14890, nc14891, nc14892, 
        nc14893, nc14894, \A_DOUT_TEMPR61[39] , \A_DOUT_TEMPR61[38] , 
        \A_DOUT_TEMPR61[37] , \A_DOUT_TEMPR61[36] , 
        \A_DOUT_TEMPR61[35] }), .B_DOUT({nc14895, nc14896, nc14897, 
        nc14898, nc14899, nc14900, nc14901, nc14902, nc14903, nc14904, 
        nc14905, nc14906, nc14907, nc14908, nc14909, 
        \B_DOUT_TEMPR61[39] , \B_DOUT_TEMPR61[38] , 
        \B_DOUT_TEMPR61[37] , \B_DOUT_TEMPR61[36] , 
        \B_DOUT_TEMPR61[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[61][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2672 (.A(\A_DOUT_TEMPR64[12] ), .B(\A_DOUT_TEMPR65[12] ), 
        .C(\A_DOUT_TEMPR66[12] ), .D(\A_DOUT_TEMPR67[12] ), .Y(
        OR4_2672_Y));
    OR4 OR4_1839 (.A(\B_DOUT_TEMPR91[2] ), .B(\B_DOUT_TEMPR92[2] ), .C(
        \B_DOUT_TEMPR93[2] ), .D(\B_DOUT_TEMPR94[2] ), .Y(OR4_1839_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%59%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R59C6 (
        .A_DOUT({nc14910, nc14911, nc14912, nc14913, nc14914, nc14915, 
        nc14916, nc14917, nc14918, nc14919, nc14920, nc14921, nc14922, 
        nc14923, nc14924, \A_DOUT_TEMPR59[34] , \A_DOUT_TEMPR59[33] , 
        \A_DOUT_TEMPR59[32] , \A_DOUT_TEMPR59[31] , 
        \A_DOUT_TEMPR59[30] }), .B_DOUT({nc14925, nc14926, nc14927, 
        nc14928, nc14929, nc14930, nc14931, nc14932, nc14933, nc14934, 
        nc14935, nc14936, nc14937, nc14938, nc14939, 
        \B_DOUT_TEMPR59[34] , \B_DOUT_TEMPR59[33] , 
        \B_DOUT_TEMPR59[32] , \B_DOUT_TEMPR59[31] , 
        \B_DOUT_TEMPR59[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[59][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1625 (.A(\A_DOUT_TEMPR68[10] ), .B(\A_DOUT_TEMPR69[10] ), 
        .C(\A_DOUT_TEMPR70[10] ), .D(\A_DOUT_TEMPR71[10] ), .Y(
        OR4_1625_Y));
    OR4 OR4_730 (.A(\A_DOUT_TEMPR8[11] ), .B(\A_DOUT_TEMPR9[11] ), .C(
        \A_DOUT_TEMPR10[11] ), .D(\A_DOUT_TEMPR11[11] ), .Y(OR4_730_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%110%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R110C6 (
        .A_DOUT({nc14940, nc14941, nc14942, nc14943, nc14944, nc14945, 
        nc14946, nc14947, nc14948, nc14949, nc14950, nc14951, nc14952, 
        nc14953, nc14954, \A_DOUT_TEMPR110[34] , \A_DOUT_TEMPR110[33] , 
        \A_DOUT_TEMPR110[32] , \A_DOUT_TEMPR110[31] , 
        \A_DOUT_TEMPR110[30] }), .B_DOUT({nc14955, nc14956, nc14957, 
        nc14958, nc14959, nc14960, nc14961, nc14962, nc14963, nc14964, 
        nc14965, nc14966, nc14967, nc14968, nc14969, 
        \B_DOUT_TEMPR110[34] , \B_DOUT_TEMPR110[33] , 
        \B_DOUT_TEMPR110[32] , \B_DOUT_TEMPR110[31] , 
        \B_DOUT_TEMPR110[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[110][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%112%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R112C6 (
        .A_DOUT({nc14970, nc14971, nc14972, nc14973, nc14974, nc14975, 
        nc14976, nc14977, nc14978, nc14979, nc14980, nc14981, nc14982, 
        nc14983, nc14984, \A_DOUT_TEMPR112[34] , \A_DOUT_TEMPR112[33] , 
        \A_DOUT_TEMPR112[32] , \A_DOUT_TEMPR112[31] , 
        \A_DOUT_TEMPR112[30] }), .B_DOUT({nc14985, nc14986, nc14987, 
        nc14988, nc14989, nc14990, nc14991, nc14992, nc14993, nc14994, 
        nc14995, nc14996, nc14997, nc14998, nc14999, 
        \B_DOUT_TEMPR112[34] , \B_DOUT_TEMPR112[33] , 
        \B_DOUT_TEMPR112[32] , \B_DOUT_TEMPR112[31] , 
        \B_DOUT_TEMPR112[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[112][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_50 (.A(\B_DOUT_TEMPR72[27] ), .B(\B_DOUT_TEMPR73[27] ), .Y(
        OR2_50_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%16%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R16C2 (
        .A_DOUT({nc15000, nc15001, nc15002, nc15003, nc15004, nc15005, 
        nc15006, nc15007, nc15008, nc15009, nc15010, nc15011, nc15012, 
        nc15013, nc15014, \A_DOUT_TEMPR16[14] , \A_DOUT_TEMPR16[13] , 
        \A_DOUT_TEMPR16[12] , \A_DOUT_TEMPR16[11] , 
        \A_DOUT_TEMPR16[10] }), .B_DOUT({nc15015, nc15016, nc15017, 
        nc15018, nc15019, nc15020, nc15021, nc15022, nc15023, nc15024, 
        nc15025, nc15026, nc15027, nc15028, nc15029, 
        \B_DOUT_TEMPR16[14] , \B_DOUT_TEMPR16[13] , 
        \B_DOUT_TEMPR16[12] , \B_DOUT_TEMPR16[11] , 
        \B_DOUT_TEMPR16[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_840 (.A(\B_DOUT_TEMPR111[20] ), .B(\B_DOUT_TEMPR112[20] ), 
        .C(\B_DOUT_TEMPR113[20] ), .D(\B_DOUT_TEMPR114[20] ), .Y(
        OR4_840_Y));
    OR4 OR4_526 (.A(\B_DOUT_TEMPR115[12] ), .B(\B_DOUT_TEMPR116[12] ), 
        .C(\B_DOUT_TEMPR117[12] ), .D(\B_DOUT_TEMPR118[12] ), .Y(
        OR4_526_Y));
    OR4 OR4_2972 (.A(\B_DOUT_TEMPR48[38] ), .B(\B_DOUT_TEMPR49[38] ), 
        .C(\B_DOUT_TEMPR50[38] ), .D(\B_DOUT_TEMPR51[38] ), .Y(
        OR4_2972_Y));
    OR4 OR4_2131 (.A(OR4_695_Y), .B(OR4_500_Y), .C(OR4_1375_Y), .D(
        OR4_2553_Y), .Y(OR4_2131_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%45%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R45C5 (
        .A_DOUT({nc15030, nc15031, nc15032, nc15033, nc15034, nc15035, 
        nc15036, nc15037, nc15038, nc15039, nc15040, nc15041, nc15042, 
        nc15043, nc15044, \A_DOUT_TEMPR45[29] , \A_DOUT_TEMPR45[28] , 
        \A_DOUT_TEMPR45[27] , \A_DOUT_TEMPR45[26] , 
        \A_DOUT_TEMPR45[25] }), .B_DOUT({nc15045, nc15046, nc15047, 
        nc15048, nc15049, nc15050, nc15051, nc15052, nc15053, nc15054, 
        nc15055, nc15056, nc15057, nc15058, nc15059, 
        \B_DOUT_TEMPR45[29] , \B_DOUT_TEMPR45[28] , 
        \B_DOUT_TEMPR45[27] , \B_DOUT_TEMPR45[26] , 
        \B_DOUT_TEMPR45[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%10%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R10C6 (
        .A_DOUT({nc15060, nc15061, nc15062, nc15063, nc15064, nc15065, 
        nc15066, nc15067, nc15068, nc15069, nc15070, nc15071, nc15072, 
        nc15073, nc15074, \A_DOUT_TEMPR10[34] , \A_DOUT_TEMPR10[33] , 
        \A_DOUT_TEMPR10[32] , \A_DOUT_TEMPR10[31] , 
        \A_DOUT_TEMPR10[30] }), .B_DOUT({nc15075, nc15076, nc15077, 
        nc15078, nc15079, nc15080, nc15081, nc15082, nc15083, nc15084, 
        nc15085, nc15086, nc15087, nc15088, nc15089, 
        \B_DOUT_TEMPR10[34] , \B_DOUT_TEMPR10[33] , 
        \B_DOUT_TEMPR10[32] , \B_DOUT_TEMPR10[31] , 
        \B_DOUT_TEMPR10[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_540 (.A(\B_DOUT_TEMPR48[22] ), .B(\B_DOUT_TEMPR49[22] ), 
        .C(\B_DOUT_TEMPR50[22] ), .D(\B_DOUT_TEMPR51[22] ), .Y(
        OR4_540_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%10%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R10C5 (
        .A_DOUT({nc15090, nc15091, nc15092, nc15093, nc15094, nc15095, 
        nc15096, nc15097, nc15098, nc15099, nc15100, nc15101, nc15102, 
        nc15103, nc15104, \A_DOUT_TEMPR10[29] , \A_DOUT_TEMPR10[28] , 
        \A_DOUT_TEMPR10[27] , \A_DOUT_TEMPR10[26] , 
        \A_DOUT_TEMPR10[25] }), .B_DOUT({nc15105, nc15106, nc15107, 
        nc15108, nc15109, nc15110, nc15111, nc15112, nc15113, nc15114, 
        nc15115, nc15116, nc15117, nc15118, nc15119, 
        \B_DOUT_TEMPR10[29] , \B_DOUT_TEMPR10[28] , 
        \B_DOUT_TEMPR10[27] , \B_DOUT_TEMPR10[26] , 
        \B_DOUT_TEMPR10[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_984 (.A(\A_DOUT_TEMPR52[21] ), .B(\A_DOUT_TEMPR53[21] ), 
        .C(\A_DOUT_TEMPR54[21] ), .D(\A_DOUT_TEMPR55[21] ), .Y(
        OR4_984_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%44%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R44C5 (
        .A_DOUT({nc15120, nc15121, nc15122, nc15123, nc15124, nc15125, 
        nc15126, nc15127, nc15128, nc15129, nc15130, nc15131, nc15132, 
        nc15133, nc15134, \A_DOUT_TEMPR44[29] , \A_DOUT_TEMPR44[28] , 
        \A_DOUT_TEMPR44[27] , \A_DOUT_TEMPR44[26] , 
        \A_DOUT_TEMPR44[25] }), .B_DOUT({nc15135, nc15136, nc15137, 
        nc15138, nc15139, nc15140, nc15141, nc15142, nc15143, nc15144, 
        nc15145, nc15146, nc15147, nc15148, nc15149, 
        \B_DOUT_TEMPR44[29] , \B_DOUT_TEMPR44[28] , 
        \B_DOUT_TEMPR44[27] , \B_DOUT_TEMPR44[26] , 
        \B_DOUT_TEMPR44[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[44][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2981 (.A(\A_DOUT_TEMPR111[8] ), .B(\A_DOUT_TEMPR112[8] ), 
        .C(\A_DOUT_TEMPR113[8] ), .D(\A_DOUT_TEMPR114[8] ), .Y(
        OR4_2981_Y));
    OR4 OR4_1131 (.A(\A_DOUT_TEMPR79[29] ), .B(\A_DOUT_TEMPR80[29] ), 
        .C(\A_DOUT_TEMPR81[29] ), .D(\A_DOUT_TEMPR82[29] ), .Y(
        OR4_1131_Y));
    OR4 OR4_2035 (.A(\A_DOUT_TEMPR12[18] ), .B(\A_DOUT_TEMPR13[18] ), 
        .C(\A_DOUT_TEMPR14[18] ), .D(\A_DOUT_TEMPR15[18] ), .Y(
        OR4_2035_Y));
    OR4 OR4_1652 (.A(\B_DOUT_TEMPR32[16] ), .B(\B_DOUT_TEMPR33[16] ), 
        .C(\B_DOUT_TEMPR34[16] ), .D(\B_DOUT_TEMPR35[16] ), .Y(
        OR4_1652_Y));
    OR4 OR4_3015 (.A(\B_DOUT_TEMPR32[37] ), .B(\B_DOUT_TEMPR33[37] ), 
        .C(\B_DOUT_TEMPR34[37] ), .D(\B_DOUT_TEMPR35[37] ), .Y(
        OR4_3015_Y));
    OR4 OR4_2293 (.A(OR4_2735_Y), .B(OR4_620_Y), .C(OR4_1115_Y), .D(
        OR4_1842_Y), .Y(OR4_2293_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%100%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R100C2 (
        .A_DOUT({nc15150, nc15151, nc15152, nc15153, nc15154, nc15155, 
        nc15156, nc15157, nc15158, nc15159, nc15160, nc15161, nc15162, 
        nc15163, nc15164, \A_DOUT_TEMPR100[14] , \A_DOUT_TEMPR100[13] , 
        \A_DOUT_TEMPR100[12] , \A_DOUT_TEMPR100[11] , 
        \A_DOUT_TEMPR100[10] }), .B_DOUT({nc15165, nc15166, nc15167, 
        nc15168, nc15169, nc15170, nc15171, nc15172, nc15173, nc15174, 
        nc15175, nc15176, nc15177, nc15178, nc15179, 
        \B_DOUT_TEMPR100[14] , \B_DOUT_TEMPR100[13] , 
        \B_DOUT_TEMPR100[12] , \B_DOUT_TEMPR100[11] , 
        \B_DOUT_TEMPR100[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[100][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_744 (.A(OR4_502_Y), .B(OR4_2063_Y), .C(OR4_2919_Y), .D(
        OR4_1914_Y), .Y(OR4_744_Y));
    OR4 OR4_1627 (.A(\B_DOUT_TEMPR40[9] ), .B(\B_DOUT_TEMPR41[9] ), .C(
        \B_DOUT_TEMPR42[9] ), .D(\B_DOUT_TEMPR43[9] ), .Y(OR4_1627_Y));
    OR4 OR4_1035 (.A(OR4_1432_Y), .B(OR4_2342_Y), .C(OR4_2001_Y), .D(
        OR4_457_Y), .Y(OR4_1035_Y));
    OR4 OR4_602 (.A(\A_DOUT_TEMPR111[24] ), .B(\A_DOUT_TEMPR112[24] ), 
        .C(\A_DOUT_TEMPR113[24] ), .D(\A_DOUT_TEMPR114[24] ), .Y(
        OR4_602_Y));
    OR4 OR4_1952 (.A(\B_DOUT_TEMPR99[3] ), .B(\B_DOUT_TEMPR100[3] ), 
        .C(\B_DOUT_TEMPR101[3] ), .D(\B_DOUT_TEMPR102[3] ), .Y(
        OR4_1952_Y));
    OR4 OR4_1107 (.A(OR4_577_Y), .B(OR4_1566_Y), .C(OR4_2223_Y), .D(
        OR4_890_Y), .Y(OR4_1107_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%110%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R110C5 (
        .A_DOUT({nc15180, nc15181, nc15182, nc15183, nc15184, nc15185, 
        nc15186, nc15187, nc15188, nc15189, nc15190, nc15191, nc15192, 
        nc15193, nc15194, \A_DOUT_TEMPR110[29] , \A_DOUT_TEMPR110[28] , 
        \A_DOUT_TEMPR110[27] , \A_DOUT_TEMPR110[26] , 
        \A_DOUT_TEMPR110[25] }), .B_DOUT({nc15195, nc15196, nc15197, 
        nc15198, nc15199, nc15200, nc15201, nc15202, nc15203, nc15204, 
        nc15205, nc15206, nc15207, nc15208, nc15209, 
        \B_DOUT_TEMPR110[29] , \B_DOUT_TEMPR110[28] , 
        \B_DOUT_TEMPR110[27] , \B_DOUT_TEMPR110[26] , 
        \B_DOUT_TEMPR110[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[110][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1604 (.A(\A_DOUT_TEMPR99[0] ), .B(\A_DOUT_TEMPR100[0] ), 
        .C(\A_DOUT_TEMPR101[0] ), .D(\A_DOUT_TEMPR102[0] ), .Y(
        OR4_1604_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%91%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R91C0 (
        .A_DOUT({nc15210, nc15211, nc15212, nc15213, nc15214, nc15215, 
        nc15216, nc15217, nc15218, nc15219, nc15220, nc15221, nc15222, 
        nc15223, nc15224, \A_DOUT_TEMPR91[4] , \A_DOUT_TEMPR91[3] , 
        \A_DOUT_TEMPR91[2] , \A_DOUT_TEMPR91[1] , \A_DOUT_TEMPR91[0] })
        , .B_DOUT({nc15225, nc15226, nc15227, nc15228, nc15229, 
        nc15230, nc15231, nc15232, nc15233, nc15234, nc15235, nc15236, 
        nc15237, nc15238, nc15239, \B_DOUT_TEMPR91[4] , 
        \B_DOUT_TEMPR91[3] , \B_DOUT_TEMPR91[2] , \B_DOUT_TEMPR91[1] , 
        \B_DOUT_TEMPR91[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[91][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_55 (.A(OR4_2114_Y), .B(OR4_66_Y), .C(OR4_743_Y), .D(
        OR4_2402_Y), .Y(OR4_55_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%57%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R57C1 (
        .A_DOUT({nc15240, nc15241, nc15242, nc15243, nc15244, nc15245, 
        nc15246, nc15247, nc15248, nc15249, nc15250, nc15251, nc15252, 
        nc15253, nc15254, \A_DOUT_TEMPR57[9] , \A_DOUT_TEMPR57[8] , 
        \A_DOUT_TEMPR57[7] , \A_DOUT_TEMPR57[6] , \A_DOUT_TEMPR57[5] })
        , .B_DOUT({nc15255, nc15256, nc15257, nc15258, nc15259, 
        nc15260, nc15261, nc15262, nc15263, nc15264, nc15265, nc15266, 
        nc15267, nc15268, nc15269, \B_DOUT_TEMPR57[9] , 
        \B_DOUT_TEMPR57[8] , \B_DOUT_TEMPR57[7] , \B_DOUT_TEMPR57[6] , 
        \B_DOUT_TEMPR57[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[57][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2837 (.A(OR4_3025_Y), .B(OR4_2839_Y), .C(OR4_649_Y), .D(
        OR4_1833_Y), .Y(OR4_2837_Y));
    OR4 OR4_2218 (.A(\A_DOUT_TEMPR95[29] ), .B(\A_DOUT_TEMPR96[29] ), 
        .C(\A_DOUT_TEMPR97[29] ), .D(\A_DOUT_TEMPR98[29] ), .Y(
        OR4_2218_Y));
    OR4 OR4_519 (.A(OR4_1311_Y), .B(OR4_2189_Y), .C(OR4_1861_Y), .D(
        OR4_304_Y), .Y(OR4_519_Y));
    OR4 OR4_1189 (.A(OR4_2905_Y), .B(OR4_2711_Y), .C(OR2_67_Y), .D(
        \B_DOUT_TEMPR74[33] ), .Y(OR4_1189_Y));
    OR4 OR4_2283 (.A(\B_DOUT_TEMPR0[21] ), .B(\B_DOUT_TEMPR1[21] ), .C(
        \B_DOUT_TEMPR2[21] ), .D(\B_DOUT_TEMPR3[21] ), .Y(OR4_2283_Y));
    OR4 OR4_1837 (.A(\B_DOUT_TEMPR52[29] ), .B(\B_DOUT_TEMPR53[29] ), 
        .C(\B_DOUT_TEMPR54[29] ), .D(\B_DOUT_TEMPR55[29] ), .Y(
        OR4_1837_Y));
    OR4 OR4_947 (.A(\B_DOUT_TEMPR99[28] ), .B(\B_DOUT_TEMPR100[28] ), 
        .C(\B_DOUT_TEMPR101[28] ), .D(\B_DOUT_TEMPR102[28] ), .Y(
        OR4_947_Y));
    OR4 OR4_2206 (.A(OR4_351_Y), .B(OR4_1670_Y), .C(OR4_1338_Y), .D(
        OR4_2363_Y), .Y(OR4_2206_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%2%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R2C1 (
        .A_DOUT({nc15270, nc15271, nc15272, nc15273, nc15274, nc15275, 
        nc15276, nc15277, nc15278, nc15279, nc15280, nc15281, nc15282, 
        nc15283, nc15284, \A_DOUT_TEMPR2[9] , \A_DOUT_TEMPR2[8] , 
        \A_DOUT_TEMPR2[7] , \A_DOUT_TEMPR2[6] , \A_DOUT_TEMPR2[5] }), 
        .B_DOUT({nc15285, nc15286, nc15287, nc15288, nc15289, nc15290, 
        nc15291, nc15292, nc15293, nc15294, nc15295, nc15296, nc15297, 
        nc15298, nc15299, \B_DOUT_TEMPR2[9] , \B_DOUT_TEMPR2[8] , 
        \B_DOUT_TEMPR2[7] , \B_DOUT_TEMPR2[6] , \B_DOUT_TEMPR2[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[2][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[0] , A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[0] , B_ADDR[13], \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1971 (.A(OR4_2550_Y), .B(OR4_2572_Y), .C(OR4_144_Y), .D(
        OR4_2372_Y), .Y(OR4_1971_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%39%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R39C6 (
        .A_DOUT({nc15300, nc15301, nc15302, nc15303, nc15304, nc15305, 
        nc15306, nc15307, nc15308, nc15309, nc15310, nc15311, nc15312, 
        nc15313, nc15314, \A_DOUT_TEMPR39[34] , \A_DOUT_TEMPR39[33] , 
        \A_DOUT_TEMPR39[32] , \A_DOUT_TEMPR39[31] , 
        \A_DOUT_TEMPR39[30] }), .B_DOUT({nc15315, nc15316, nc15317, 
        nc15318, nc15319, nc15320, nc15321, nc15322, nc15323, nc15324, 
        nc15325, nc15326, nc15327, nc15328, nc15329, 
        \B_DOUT_TEMPR39[34] , \B_DOUT_TEMPR39[33] , 
        \B_DOUT_TEMPR39[32] , \B_DOUT_TEMPR39[31] , 
        \B_DOUT_TEMPR39[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[39][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%115%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R115C2 (
        .A_DOUT({nc15330, nc15331, nc15332, nc15333, nc15334, nc15335, 
        nc15336, nc15337, nc15338, nc15339, nc15340, nc15341, nc15342, 
        nc15343, nc15344, \A_DOUT_TEMPR115[14] , \A_DOUT_TEMPR115[13] , 
        \A_DOUT_TEMPR115[12] , \A_DOUT_TEMPR115[11] , 
        \A_DOUT_TEMPR115[10] }), .B_DOUT({nc15345, nc15346, nc15347, 
        nc15348, nc15349, nc15350, nc15351, nc15352, nc15353, nc15354, 
        nc15355, nc15356, nc15357, nc15358, nc15359, 
        \B_DOUT_TEMPR115[14] , \B_DOUT_TEMPR115[13] , 
        \B_DOUT_TEMPR115[12] , \B_DOUT_TEMPR115[11] , 
        \B_DOUT_TEMPR115[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[115][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2544 (.A(\B_DOUT_TEMPR24[31] ), .B(\B_DOUT_TEMPR25[31] ), 
        .C(\B_DOUT_TEMPR26[31] ), .D(\B_DOUT_TEMPR27[31] ), .Y(
        OR4_2544_Y));
    OR4 OR4_1993 (.A(OR4_865_Y), .B(OR4_47_Y), .C(OR4_2048_Y), .D(
        OR4_2343_Y), .Y(OR4_1993_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%118%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R118C0 (
        .A_DOUT({nc15360, nc15361, nc15362, nc15363, nc15364, nc15365, 
        nc15366, nc15367, nc15368, nc15369, nc15370, nc15371, nc15372, 
        nc15373, nc15374, \A_DOUT_TEMPR118[4] , \A_DOUT_TEMPR118[3] , 
        \A_DOUT_TEMPR118[2] , \A_DOUT_TEMPR118[1] , 
        \A_DOUT_TEMPR118[0] }), .B_DOUT({nc15375, nc15376, nc15377, 
        nc15378, nc15379, nc15380, nc15381, nc15382, nc15383, nc15384, 
        nc15385, nc15386, nc15387, nc15388, nc15389, 
        \B_DOUT_TEMPR118[4] , \B_DOUT_TEMPR118[3] , 
        \B_DOUT_TEMPR118[2] , \B_DOUT_TEMPR118[1] , 
        \B_DOUT_TEMPR118[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[118][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%67%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R67C0 (
        .A_DOUT({nc15390, nc15391, nc15392, nc15393, nc15394, nc15395, 
        nc15396, nc15397, nc15398, nc15399, nc15400, nc15401, nc15402, 
        nc15403, nc15404, \A_DOUT_TEMPR67[4] , \A_DOUT_TEMPR67[3] , 
        \A_DOUT_TEMPR67[2] , \A_DOUT_TEMPR67[1] , \A_DOUT_TEMPR67[0] })
        , .B_DOUT({nc15405, nc15406, nc15407, nc15408, nc15409, 
        nc15410, nc15411, nc15412, nc15413, nc15414, nc15415, nc15416, 
        nc15417, nc15418, nc15419, \B_DOUT_TEMPR67[4] , 
        \B_DOUT_TEMPR67[3] , \B_DOUT_TEMPR67[2] , \B_DOUT_TEMPR67[1] , 
        \B_DOUT_TEMPR67[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[67][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_546 (.A(\A_DOUT_TEMPR40[32] ), .B(\A_DOUT_TEMPR41[32] ), 
        .C(\A_DOUT_TEMPR42[32] ), .D(\A_DOUT_TEMPR43[32] ), .Y(
        OR4_546_Y));
    OR4 OR4_2479 (.A(\B_DOUT_TEMPR16[5] ), .B(\B_DOUT_TEMPR17[5] ), .C(
        \B_DOUT_TEMPR18[5] ), .D(\B_DOUT_TEMPR19[5] ), .Y(OR4_2479_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%18%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R18C5 (
        .A_DOUT({nc15420, nc15421, nc15422, nc15423, nc15424, nc15425, 
        nc15426, nc15427, nc15428, nc15429, nc15430, nc15431, nc15432, 
        nc15433, nc15434, \A_DOUT_TEMPR18[29] , \A_DOUT_TEMPR18[28] , 
        \A_DOUT_TEMPR18[27] , \A_DOUT_TEMPR18[26] , 
        \A_DOUT_TEMPR18[25] }), .B_DOUT({nc15435, nc15436, nc15437, 
        nc15438, nc15439, nc15440, nc15441, nc15442, nc15443, nc15444, 
        nc15445, nc15446, nc15447, nc15448, nc15449, 
        \B_DOUT_TEMPR18[29] , \B_DOUT_TEMPR18[28] , 
        \B_DOUT_TEMPR18[27] , \B_DOUT_TEMPR18[26] , 
        \B_DOUT_TEMPR18[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_78 (.A(\B_DOUT_TEMPR72[3] ), .B(\B_DOUT_TEMPR73[3] ), .Y(
        OR2_78_Y));
    OR4 OR4_1391 (.A(\B_DOUT_TEMPR40[15] ), .B(\B_DOUT_TEMPR41[15] ), 
        .C(\B_DOUT_TEMPR42[15] ), .D(\B_DOUT_TEMPR43[15] ), .Y(
        OR4_1391_Y));
    OR4 OR4_1324 (.A(\B_DOUT_TEMPR28[11] ), .B(\B_DOUT_TEMPR29[11] ), 
        .C(\B_DOUT_TEMPR30[11] ), .D(\B_DOUT_TEMPR31[11] ), .Y(
        OR4_1324_Y));
    OR4 OR4_2129 (.A(\B_DOUT_TEMPR32[0] ), .B(\B_DOUT_TEMPR33[0] ), .C(
        \B_DOUT_TEMPR34[0] ), .D(\B_DOUT_TEMPR35[0] ), .Y(OR4_2129_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%48%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R48C4 (
        .A_DOUT({nc15450, nc15451, nc15452, nc15453, nc15454, nc15455, 
        nc15456, nc15457, nc15458, nc15459, nc15460, nc15461, nc15462, 
        nc15463, nc15464, \A_DOUT_TEMPR48[24] , \A_DOUT_TEMPR48[23] , 
        \A_DOUT_TEMPR48[22] , \A_DOUT_TEMPR48[21] , 
        \A_DOUT_TEMPR48[20] }), .B_DOUT({nc15465, nc15466, nc15467, 
        nc15468, nc15469, nc15470, nc15471, nc15472, nc15473, nc15474, 
        nc15475, nc15476, nc15477, nc15478, nc15479, 
        \B_DOUT_TEMPR48[24] , \B_DOUT_TEMPR48[23] , 
        \B_DOUT_TEMPR48[22] , \B_DOUT_TEMPR48[21] , 
        \B_DOUT_TEMPR48[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[48][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_55 (.A(\B_DOUT_TEMPR72[16] ), .B(\B_DOUT_TEMPR73[16] ), .Y(
        OR2_55_Y));
    OR4 OR4_1273 (.A(OR4_1692_Y), .B(OR4_2090_Y), .C(OR4_2859_Y), .D(
        OR4_611_Y), .Y(OR4_1273_Y));
    OR4 OR4_1891 (.A(\A_DOUT_TEMPR40[14] ), .B(\A_DOUT_TEMPR41[14] ), 
        .C(\A_DOUT_TEMPR42[14] ), .D(\A_DOUT_TEMPR43[14] ), .Y(
        OR4_1891_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%4%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R4C5 (
        .A_DOUT({nc15480, nc15481, nc15482, nc15483, nc15484, nc15485, 
        nc15486, nc15487, nc15488, nc15489, nc15490, nc15491, nc15492, 
        nc15493, nc15494, \A_DOUT_TEMPR4[29] , \A_DOUT_TEMPR4[28] , 
        \A_DOUT_TEMPR4[27] , \A_DOUT_TEMPR4[26] , \A_DOUT_TEMPR4[25] })
        , .B_DOUT({nc15495, nc15496, nc15497, nc15498, nc15499, 
        nc15500, nc15501, nc15502, nc15503, nc15504, nc15505, nc15506, 
        nc15507, nc15508, nc15509, \B_DOUT_TEMPR4[29] , 
        \B_DOUT_TEMPR4[28] , \B_DOUT_TEMPR4[27] , \B_DOUT_TEMPR4[26] , 
        \B_DOUT_TEMPR4[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1459 (.A(\A_DOUT_TEMPR60[32] ), .B(\A_DOUT_TEMPR61[32] ), 
        .C(\A_DOUT_TEMPR62[32] ), .D(\A_DOUT_TEMPR63[32] ), .Y(
        OR4_1459_Y));
    OR4 OR4_468 (.A(\B_DOUT_TEMPR16[31] ), .B(\B_DOUT_TEMPR17[31] ), 
        .C(\B_DOUT_TEMPR18[31] ), .D(\B_DOUT_TEMPR19[31] ), .Y(
        OR4_468_Y));
    OR4 OR4_2806 (.A(OR4_539_Y), .B(OR4_2610_Y), .C(OR4_2828_Y), .D(
        OR4_2618_Y), .Y(OR4_2806_Y));
    OR4 OR4_2241 (.A(\B_DOUT_TEMPR52[16] ), .B(\B_DOUT_TEMPR53[16] ), 
        .C(\B_DOUT_TEMPR54[16] ), .D(\B_DOUT_TEMPR55[16] ), .Y(
        OR4_2241_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%7%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R7C4 (
        .A_DOUT({nc15510, nc15511, nc15512, nc15513, nc15514, nc15515, 
        nc15516, nc15517, nc15518, nc15519, nc15520, nc15521, nc15522, 
        nc15523, nc15524, \A_DOUT_TEMPR7[24] , \A_DOUT_TEMPR7[23] , 
        \A_DOUT_TEMPR7[22] , \A_DOUT_TEMPR7[21] , \A_DOUT_TEMPR7[20] })
        , .B_DOUT({nc15525, nc15526, nc15527, nc15528, nc15529, 
        nc15530, nc15531, nc15532, nc15533, nc15534, nc15535, nc15536, 
        nc15537, nc15538, nc15539, \B_DOUT_TEMPR7[24] , 
        \B_DOUT_TEMPR7[23] , \B_DOUT_TEMPR7[22] , \B_DOUT_TEMPR7[21] , 
        \B_DOUT_TEMPR7[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_564 (.A(\B_DOUT_TEMPR87[12] ), .B(\B_DOUT_TEMPR88[12] ), 
        .C(\B_DOUT_TEMPR89[12] ), .D(\B_DOUT_TEMPR90[12] ), .Y(
        OR4_564_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%37%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R37C1 (
        .A_DOUT({nc15540, nc15541, nc15542, nc15543, nc15544, nc15545, 
        nc15546, nc15547, nc15548, nc15549, nc15550, nc15551, nc15552, 
        nc15553, nc15554, \A_DOUT_TEMPR37[9] , \A_DOUT_TEMPR37[8] , 
        \A_DOUT_TEMPR37[7] , \A_DOUT_TEMPR37[6] , \A_DOUT_TEMPR37[5] })
        , .B_DOUT({nc15555, nc15556, nc15557, nc15558, nc15559, 
        nc15560, nc15561, nc15562, nc15563, nc15564, nc15565, nc15566, 
        nc15567, nc15568, nc15569, \B_DOUT_TEMPR37[9] , 
        \B_DOUT_TEMPR37[8] , \B_DOUT_TEMPR37[7] , \B_DOUT_TEMPR37[6] , 
        \B_DOUT_TEMPR37[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[37][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2370 (.A(\B_DOUT_TEMPR87[30] ), .B(\B_DOUT_TEMPR88[30] ), 
        .C(\B_DOUT_TEMPR89[30] ), .D(\B_DOUT_TEMPR90[30] ), .Y(
        OR4_2370_Y));
    OR4 OR4_2477 (.A(\B_DOUT_TEMPR4[32] ), .B(\B_DOUT_TEMPR5[32] ), .C(
        \B_DOUT_TEMPR6[32] ), .D(\B_DOUT_TEMPR7[32] ), .Y(OR4_2477_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%11%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R11C7 (
        .A_DOUT({nc15570, nc15571, nc15572, nc15573, nc15574, nc15575, 
        nc15576, nc15577, nc15578, nc15579, nc15580, nc15581, nc15582, 
        nc15583, nc15584, \A_DOUT_TEMPR11[39] , \A_DOUT_TEMPR11[38] , 
        \A_DOUT_TEMPR11[37] , \A_DOUT_TEMPR11[36] , 
        \A_DOUT_TEMPR11[35] }), .B_DOUT({nc15585, nc15586, nc15587, 
        nc15588, nc15589, nc15590, nc15591, nc15592, nc15593, nc15594, 
        nc15595, nc15596, nc15597, nc15598, nc15599, 
        \B_DOUT_TEMPR11[39] , \B_DOUT_TEMPR11[38] , 
        \B_DOUT_TEMPR11[37] , \B_DOUT_TEMPR11[36] , 
        \B_DOUT_TEMPR11[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[39]  (.A(OR4_2527_Y), .B(OR4_2187_Y), .C(
        OR4_2069_Y), .D(OR4_1200_Y), .Y(A_DOUT[39]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%84%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R84C0 (
        .A_DOUT({nc15600, nc15601, nc15602, nc15603, nc15604, nc15605, 
        nc15606, nc15607, nc15608, nc15609, nc15610, nc15611, nc15612, 
        nc15613, nc15614, \A_DOUT_TEMPR84[4] , \A_DOUT_TEMPR84[3] , 
        \A_DOUT_TEMPR84[2] , \A_DOUT_TEMPR84[1] , \A_DOUT_TEMPR84[0] })
        , .B_DOUT({nc15615, nc15616, nc15617, nc15618, nc15619, 
        nc15620, nc15621, nc15622, nc15623, nc15624, nc15625, nc15626, 
        nc15627, nc15628, nc15629, \B_DOUT_TEMPR84[4] , 
        \B_DOUT_TEMPR84[3] , \B_DOUT_TEMPR84[2] , \B_DOUT_TEMPR84[1] , 
        \B_DOUT_TEMPR84[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[84][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%117%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R117C6 (
        .A_DOUT({nc15630, nc15631, nc15632, nc15633, nc15634, nc15635, 
        nc15636, nc15637, nc15638, nc15639, nc15640, nc15641, nc15642, 
        nc15643, nc15644, \A_DOUT_TEMPR117[34] , \A_DOUT_TEMPR117[33] , 
        \A_DOUT_TEMPR117[32] , \A_DOUT_TEMPR117[31] , 
        \A_DOUT_TEMPR117[30] }), .B_DOUT({nc15645, nc15646, nc15647, 
        nc15648, nc15649, nc15650, nc15651, nc15652, nc15653, nc15654, 
        nc15655, nc15656, nc15657, nc15658, nc15659, 
        \B_DOUT_TEMPR117[34] , \B_DOUT_TEMPR117[33] , 
        \B_DOUT_TEMPR117[32] , \B_DOUT_TEMPR117[31] , 
        \B_DOUT_TEMPR117[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[117][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_652 (.A(OR4_2932_Y), .B(OR4_839_Y), .C(OR4_114_Y), .D(
        OR4_2880_Y), .Y(OR4_652_Y));
    OR2 OR2_31 (.A(\A_DOUT_TEMPR72[23] ), .B(\A_DOUT_TEMPR73[23] ), .Y(
        OR2_31_Y));
    OR4 OR4_1168 (.A(\A_DOUT_TEMPR107[29] ), .B(\A_DOUT_TEMPR108[29] ), 
        .C(\A_DOUT_TEMPR109[29] ), .D(\A_DOUT_TEMPR110[29] ), .Y(
        OR4_1168_Y));
    OR4 OR4_1019 (.A(\B_DOUT_TEMPR56[35] ), .B(\B_DOUT_TEMPR57[35] ), 
        .C(\B_DOUT_TEMPR58[35] ), .D(\B_DOUT_TEMPR59[35] ), .Y(
        OR4_1019_Y));
    OR4 OR4_1350 (.A(\A_DOUT_TEMPR79[35] ), .B(\A_DOUT_TEMPR80[35] ), 
        .C(\A_DOUT_TEMPR81[35] ), .D(\A_DOUT_TEMPR82[35] ), .Y(
        OR4_1350_Y));
    OR4 OR4_1457 (.A(\B_DOUT_TEMPR99[35] ), .B(\B_DOUT_TEMPR100[35] ), 
        .C(\B_DOUT_TEMPR101[35] ), .D(\B_DOUT_TEMPR102[35] ), .Y(
        OR4_1457_Y));
    OR4 OR4_1882 (.A(\B_DOUT_TEMPR75[33] ), .B(\B_DOUT_TEMPR76[33] ), 
        .C(\B_DOUT_TEMPR77[33] ), .D(\B_DOUT_TEMPR78[33] ), .Y(
        OR4_1882_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%73%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R73C5 (
        .A_DOUT({nc15660, nc15661, nc15662, nc15663, nc15664, nc15665, 
        nc15666, nc15667, nc15668, nc15669, nc15670, nc15671, nc15672, 
        nc15673, nc15674, \A_DOUT_TEMPR73[29] , \A_DOUT_TEMPR73[28] , 
        \A_DOUT_TEMPR73[27] , \A_DOUT_TEMPR73[26] , 
        \A_DOUT_TEMPR73[25] }), .B_DOUT({nc15675, nc15676, nc15677, 
        nc15678, nc15679, nc15680, nc15681, nc15682, nc15683, nc15684, 
        nc15685, nc15686, nc15687, nc15688, nc15689, 
        \B_DOUT_TEMPR73[29] , \B_DOUT_TEMPR73[28] , 
        \B_DOUT_TEMPR73[27] , \B_DOUT_TEMPR73[26] , 
        \B_DOUT_TEMPR73[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[73][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1600 (.A(\A_DOUT_TEMPR48[19] ), .B(\A_DOUT_TEMPR49[19] ), 
        .C(\A_DOUT_TEMPR50[19] ), .D(\A_DOUT_TEMPR51[19] ), .Y(
        OR4_1600_Y));
    OR4 OR4_489 (.A(\A_DOUT_TEMPR103[26] ), .B(\A_DOUT_TEMPR104[26] ), 
        .C(\A_DOUT_TEMPR105[26] ), .D(\A_DOUT_TEMPR106[26] ), .Y(
        OR4_489_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%86%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R86C7 (
        .A_DOUT({nc15690, nc15691, nc15692, nc15693, nc15694, nc15695, 
        nc15696, nc15697, nc15698, nc15699, nc15700, nc15701, nc15702, 
        nc15703, nc15704, \A_DOUT_TEMPR86[39] , \A_DOUT_TEMPR86[38] , 
        \A_DOUT_TEMPR86[37] , \A_DOUT_TEMPR86[36] , 
        \A_DOUT_TEMPR86[35] }), .B_DOUT({nc15705, nc15706, nc15707, 
        nc15708, nc15709, nc15710, nc15711, nc15712, nc15713, nc15714, 
        nc15715, nc15716, nc15717, nc15718, nc15719, 
        \B_DOUT_TEMPR86[39] , \B_DOUT_TEMPR86[38] , 
        \B_DOUT_TEMPR86[37] , \B_DOUT_TEMPR86[36] , 
        \B_DOUT_TEMPR86[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[86][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1519 (.A(\B_DOUT_TEMPR24[21] ), .B(\B_DOUT_TEMPR25[21] ), 
        .C(\B_DOUT_TEMPR26[21] ), .D(\B_DOUT_TEMPR27[21] ), .Y(
        OR4_1519_Y));
    OR4 OR4_2961 (.A(\B_DOUT_TEMPR36[15] ), .B(\B_DOUT_TEMPR37[15] ), 
        .C(\B_DOUT_TEMPR38[15] ), .D(\B_DOUT_TEMPR39[15] ), .Y(
        OR4_2961_Y));
    OR4 OR4_1008 (.A(\A_DOUT_TEMPR12[35] ), .B(\A_DOUT_TEMPR13[35] ), 
        .C(\A_DOUT_TEMPR14[35] ), .D(\A_DOUT_TEMPR15[35] ), .Y(
        OR4_1008_Y));
    OR4 OR4_2700 (.A(OR4_1583_Y), .B(OR4_2590_Y), .C(OR4_213_Y), .D(
        OR4_1889_Y), .Y(OR4_2700_Y));
    OR4 OR4_372 (.A(OR4_1353_Y), .B(OR4_2670_Y), .C(OR4_2290_Y), .D(
        OR4_299_Y), .Y(OR4_372_Y));
    OR4 OR4_59 (.A(\B_DOUT_TEMPR60[17] ), .B(\B_DOUT_TEMPR61[17] ), .C(
        \B_DOUT_TEMPR62[17] ), .D(\B_DOUT_TEMPR63[17] ), .Y(OR4_59_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%87%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R87C6 (
        .A_DOUT({nc15720, nc15721, nc15722, nc15723, nc15724, nc15725, 
        nc15726, nc15727, nc15728, nc15729, nc15730, nc15731, nc15732, 
        nc15733, nc15734, \A_DOUT_TEMPR87[34] , \A_DOUT_TEMPR87[33] , 
        \A_DOUT_TEMPR87[32] , \A_DOUT_TEMPR87[31] , 
        \A_DOUT_TEMPR87[30] }), .B_DOUT({nc15735, nc15736, nc15737, 
        nc15738, nc15739, nc15740, nc15741, nc15742, nc15743, nc15744, 
        nc15745, nc15746, nc15747, nc15748, nc15749, 
        \B_DOUT_TEMPR87[34] , \B_DOUT_TEMPR87[33] , 
        \B_DOUT_TEMPR87[32] , \B_DOUT_TEMPR87[31] , 
        \B_DOUT_TEMPR87[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[87][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_120 (.A(\B_DOUT_TEMPR68[37] ), .B(\B_DOUT_TEMPR69[37] ), 
        .C(\B_DOUT_TEMPR70[37] ), .D(\B_DOUT_TEMPR71[37] ), .Y(
        OR4_120_Y));
    OR4 OR4_1863 (.A(OR4_1037_Y), .B(OR4_2702_Y), .C(OR4_2121_Y), .D(
        OR4_405_Y), .Y(OR4_1863_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%44%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R44C7 (
        .A_DOUT({nc15750, nc15751, nc15752, nc15753, nc15754, nc15755, 
        nc15756, nc15757, nc15758, nc15759, nc15760, nc15761, nc15762, 
        nc15763, nc15764, \A_DOUT_TEMPR44[39] , \A_DOUT_TEMPR44[38] , 
        \A_DOUT_TEMPR44[37] , \A_DOUT_TEMPR44[36] , 
        \A_DOUT_TEMPR44[35] }), .B_DOUT({nc15765, nc15766, nc15767, 
        nc15768, nc15769, nc15770, nc15771, nc15772, nc15773, nc15774, 
        nc15775, nc15776, nc15777, nc15778, nc15779, 
        \B_DOUT_TEMPR44[39] , \B_DOUT_TEMPR44[38] , 
        \B_DOUT_TEMPR44[37] , \B_DOUT_TEMPR44[36] , 
        \B_DOUT_TEMPR44[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[44][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1312 (.A(OR4_1144_Y), .B(OR4_2170_Y), .C(OR4_2843_Y), .D(
        OR4_2008_Y), .Y(OR4_1312_Y));
    OR4 OR4_413 (.A(\B_DOUT_TEMPR99[5] ), .B(\B_DOUT_TEMPR100[5] ), .C(
        \B_DOUT_TEMPR101[5] ), .D(\B_DOUT_TEMPR102[5] ), .Y(OR4_413_Y));
    OR4 OR4_1769 (.A(\A_DOUT_TEMPR64[17] ), .B(\A_DOUT_TEMPR65[17] ), 
        .C(\A_DOUT_TEMPR66[17] ), .D(\A_DOUT_TEMPR67[17] ), .Y(
        OR4_1769_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%82%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R82C4 (
        .A_DOUT({nc15780, nc15781, nc15782, nc15783, nc15784, nc15785, 
        nc15786, nc15787, nc15788, nc15789, nc15790, nc15791, nc15792, 
        nc15793, nc15794, \A_DOUT_TEMPR82[24] , \A_DOUT_TEMPR82[23] , 
        \A_DOUT_TEMPR82[22] , \A_DOUT_TEMPR82[21] , 
        \A_DOUT_TEMPR82[20] }), .B_DOUT({nc15795, nc15796, nc15797, 
        nc15798, nc15799, nc15800, nc15801, nc15802, nc15803, nc15804, 
        nc15805, nc15806, nc15807, nc15808, nc15809, 
        \B_DOUT_TEMPR82[24] , \B_DOUT_TEMPR82[23] , 
        \B_DOUT_TEMPR82[22] , \B_DOUT_TEMPR82[21] , 
        \B_DOUT_TEMPR82[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[82][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2059 (.A(\A_DOUT_TEMPR115[17] ), .B(\A_DOUT_TEMPR116[17] ), 
        .C(\A_DOUT_TEMPR117[17] ), .D(\A_DOUT_TEMPR118[17] ), .Y(
        OR4_2059_Y));
    OR4 OR4_569 (.A(\B_DOUT_TEMPR0[28] ), .B(\B_DOUT_TEMPR1[28] ), .C(
        \B_DOUT_TEMPR2[28] ), .D(\B_DOUT_TEMPR3[28] ), .Y(OR4_569_Y));
    OR4 OR4_1683 (.A(\B_DOUT_TEMPR36[31] ), .B(\B_DOUT_TEMPR37[31] ), 
        .C(\B_DOUT_TEMPR38[31] ), .D(\B_DOUT_TEMPR39[31] ), .Y(
        OR4_1683_Y));
    OR4 OR4_181 (.A(\A_DOUT_TEMPR87[12] ), .B(\A_DOUT_TEMPR88[12] ), 
        .C(\A_DOUT_TEMPR89[12] ), .D(\A_DOUT_TEMPR90[12] ), .Y(
        OR4_181_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%76%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R76C4 (
        .A_DOUT({nc15810, nc15811, nc15812, nc15813, nc15814, nc15815, 
        nc15816, nc15817, nc15818, nc15819, nc15820, nc15821, nc15822, 
        nc15823, nc15824, \A_DOUT_TEMPR76[24] , \A_DOUT_TEMPR76[23] , 
        \A_DOUT_TEMPR76[22] , \A_DOUT_TEMPR76[21] , 
        \A_DOUT_TEMPR76[20] }), .B_DOUT({nc15825, nc15826, nc15827, 
        nc15828, nc15829, nc15830, nc15831, nc15832, nc15833, nc15834, 
        nc15835, nc15836, nc15837, nc15838, nc15839, 
        \B_DOUT_TEMPR76[24] , \B_DOUT_TEMPR76[23] , 
        \B_DOUT_TEMPR76[22] , \B_DOUT_TEMPR76[21] , 
        \B_DOUT_TEMPR76[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[76][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_628 (.A(\A_DOUT_TEMPR75[26] ), .B(\A_DOUT_TEMPR76[26] ), 
        .C(\A_DOUT_TEMPR77[26] ), .D(\A_DOUT_TEMPR78[26] ), .Y(
        OR4_628_Y));
    OR4 OR4_1420 (.A(\B_DOUT_TEMPR44[32] ), .B(\B_DOUT_TEMPR45[32] ), 
        .C(\B_DOUT_TEMPR46[32] ), .D(\B_DOUT_TEMPR47[32] ), .Y(
        OR4_1420_Y));
    OR4 OR4_2559 (.A(\B_DOUT_TEMPR8[16] ), .B(\B_DOUT_TEMPR9[16] ), .C(
        \B_DOUT_TEMPR10[16] ), .D(\B_DOUT_TEMPR11[16] ), .Y(OR4_2559_Y)
        );
    OR4 OR4_1989 (.A(\A_DOUT_TEMPR103[28] ), .B(\A_DOUT_TEMPR104[28] ), 
        .C(\A_DOUT_TEMPR105[28] ), .D(\A_DOUT_TEMPR106[28] ), .Y(
        OR4_1989_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%97%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R97C4 (
        .A_DOUT({nc15840, nc15841, nc15842, nc15843, nc15844, nc15845, 
        nc15846, nc15847, nc15848, nc15849, nc15850, nc15851, nc15852, 
        nc15853, nc15854, \A_DOUT_TEMPR97[24] , \A_DOUT_TEMPR97[23] , 
        \A_DOUT_TEMPR97[22] , \A_DOUT_TEMPR97[21] , 
        \A_DOUT_TEMPR97[20] }), .B_DOUT({nc15855, nc15856, nc15857, 
        nc15858, nc15859, nc15860, nc15861, nc15862, nc15863, nc15864, 
        nc15865, nc15866, nc15867, nc15868, nc15869, 
        \B_DOUT_TEMPR97[24] , \B_DOUT_TEMPR97[23] , 
        \B_DOUT_TEMPR97[22] , \B_DOUT_TEMPR97[21] , 
        \B_DOUT_TEMPR97[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[97][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2263 (.A(OR4_1385_Y), .B(OR4_2262_Y), .C(OR4_1454_Y), .D(
        OR4_393_Y), .Y(OR4_2263_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%69%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R69C6 (
        .A_DOUT({nc15870, nc15871, nc15872, nc15873, nc15874, nc15875, 
        nc15876, nc15877, nc15878, nc15879, nc15880, nc15881, nc15882, 
        nc15883, nc15884, \A_DOUT_TEMPR69[34] , \A_DOUT_TEMPR69[33] , 
        \A_DOUT_TEMPR69[32] , \A_DOUT_TEMPR69[31] , 
        \A_DOUT_TEMPR69[30] }), .B_DOUT({nc15885, nc15886, nc15887, 
        nc15888, nc15889, nc15890, nc15891, nc15892, nc15893, nc15894, 
        nc15895, nc15896, nc15897, nc15898, nc15899, 
        \B_DOUT_TEMPR69[34] , \B_DOUT_TEMPR69[33] , 
        \B_DOUT_TEMPR69[32] , \B_DOUT_TEMPR69[31] , 
        \B_DOUT_TEMPR69[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[69][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2822 (.A(\B_DOUT_TEMPR111[11] ), .B(\B_DOUT_TEMPR112[11] ), 
        .C(\B_DOUT_TEMPR113[11] ), .D(\B_DOUT_TEMPR114[11] ), .Y(
        OR4_2822_Y));
    OR4 OR4_1166 (.A(\A_DOUT_TEMPR36[3] ), .B(\A_DOUT_TEMPR37[3] ), .C(
        \A_DOUT_TEMPR38[3] ), .D(\A_DOUT_TEMPR39[3] ), .Y(OR4_1166_Y));
    CFG3 #( .INIT(8'h4) )  CFG3_22 (.A(B_ADDR[16]), .B(B_ADDR[15]), .C(
        B_ADDR[14]), .Y(CFG3_22_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%51%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R51C0 (
        .A_DOUT({nc15900, nc15901, nc15902, nc15903, nc15904, nc15905, 
        nc15906, nc15907, nc15908, nc15909, nc15910, nc15911, nc15912, 
        nc15913, nc15914, \A_DOUT_TEMPR51[4] , \A_DOUT_TEMPR51[3] , 
        \A_DOUT_TEMPR51[2] , \A_DOUT_TEMPR51[1] , \A_DOUT_TEMPR51[0] })
        , .B_DOUT({nc15915, nc15916, nc15917, nc15918, nc15919, 
        nc15920, nc15921, nc15922, nc15923, nc15924, nc15925, nc15926, 
        nc15927, nc15928, nc15929, \B_DOUT_TEMPR51[4] , 
        \B_DOUT_TEMPR51[3] , \B_DOUT_TEMPR51[2] , \B_DOUT_TEMPR51[1] , 
        \B_DOUT_TEMPR51[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[51][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1568 (.A(\B_DOUT_TEMPR40[35] ), .B(\B_DOUT_TEMPR41[35] ), 
        .C(\B_DOUT_TEMPR42[35] ), .D(\B_DOUT_TEMPR43[35] ), .Y(
        OR4_1568_Y));
    OR4 OR4_136 (.A(OR4_2140_Y), .B(OR4_886_Y), .C(OR4_1498_Y), .D(
        OR4_694_Y), .Y(OR4_136_Y));
    OR4 OR4_2307 (.A(OR4_1359_Y), .B(OR4_1171_Y), .C(OR4_2023_Y), .D(
        OR4_157_Y), .Y(OR4_2307_Y));
    OR4 OR4_2791 (.A(OR4_645_Y), .B(OR4_1824_Y), .C(OR2_74_Y), .D(
        \B_DOUT_TEMPR74[15] ), .Y(OR4_2791_Y));
    OR4 OR4_2202 (.A(\A_DOUT_TEMPR52[36] ), .B(\A_DOUT_TEMPR53[36] ), 
        .C(\A_DOUT_TEMPR54[36] ), .D(\A_DOUT_TEMPR55[36] ), .Y(
        OR4_2202_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%29%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R29C7 (
        .A_DOUT({nc15930, nc15931, nc15932, nc15933, nc15934, nc15935, 
        nc15936, nc15937, nc15938, nc15939, nc15940, nc15941, nc15942, 
        nc15943, nc15944, \A_DOUT_TEMPR29[39] , \A_DOUT_TEMPR29[38] , 
        \A_DOUT_TEMPR29[37] , \A_DOUT_TEMPR29[36] , 
        \A_DOUT_TEMPR29[35] }), .B_DOUT({nc15945, nc15946, nc15947, 
        nc15948, nc15949, nc15950, nc15951, nc15952, nc15953, nc15954, 
        nc15955, nc15956, nc15957, nc15958, nc15959, 
        \B_DOUT_TEMPR29[39] , \B_DOUT_TEMPR29[38] , 
        \B_DOUT_TEMPR29[37] , \B_DOUT_TEMPR29[36] , 
        \B_DOUT_TEMPR29[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_575 (.A(OR4_2439_Y), .B(OR4_674_Y), .C(OR4_1377_Y), .D(
        OR4_1653_Y), .Y(OR4_575_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%75%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R75C5 (
        .A_DOUT({nc15960, nc15961, nc15962, nc15963, nc15964, nc15965, 
        nc15966, nc15967, nc15968, nc15969, nc15970, nc15971, nc15972, 
        nc15973, nc15974, \A_DOUT_TEMPR75[29] , \A_DOUT_TEMPR75[28] , 
        \A_DOUT_TEMPR75[27] , \A_DOUT_TEMPR75[26] , 
        \A_DOUT_TEMPR75[25] }), .B_DOUT({nc15975, nc15976, nc15977, 
        nc15978, nc15979, nc15980, nc15981, nc15982, nc15983, nc15984, 
        nc15985, nc15986, nc15987, nc15988, nc15989, 
        \B_DOUT_TEMPR75[29] , \B_DOUT_TEMPR75[28] , 
        \B_DOUT_TEMPR75[27] , \B_DOUT_TEMPR75[26] , 
        \B_DOUT_TEMPR75[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[75][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%17%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R17C0 (
        .A_DOUT({nc15990, nc15991, nc15992, nc15993, nc15994, nc15995, 
        nc15996, nc15997, nc15998, nc15999, nc16000, nc16001, nc16002, 
        nc16003, nc16004, \A_DOUT_TEMPR17[4] , \A_DOUT_TEMPR17[3] , 
        \A_DOUT_TEMPR17[2] , \A_DOUT_TEMPR17[1] , \A_DOUT_TEMPR17[0] })
        , .B_DOUT({nc16005, nc16006, nc16007, nc16008, nc16009, 
        nc16010, nc16011, nc16012, nc16013, nc16014, nc16015, nc16016, 
        nc16017, nc16018, nc16019, \B_DOUT_TEMPR17[4] , 
        \B_DOUT_TEMPR17[3] , \B_DOUT_TEMPR17[2] , \B_DOUT_TEMPR17[1] , 
        \B_DOUT_TEMPR17[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h4) )  CFG3_10 (.A(A_ADDR[16]), .B(A_ADDR[15]), .C(
        A_ADDR[14]), .Y(CFG3_10_Y));
    OR4 OR4_1104 (.A(\A_DOUT_TEMPR91[19] ), .B(\A_DOUT_TEMPR92[19] ), 
        .C(\A_DOUT_TEMPR93[19] ), .D(\A_DOUT_TEMPR94[19] ), .Y(
        OR4_1104_Y));
    OR4 OR4_2352 (.A(\B_DOUT_TEMPR115[27] ), .B(\B_DOUT_TEMPR116[27] ), 
        .C(\B_DOUT_TEMPR117[27] ), .D(\B_DOUT_TEMPR118[27] ), .Y(
        OR4_2352_Y));
    OR4 OR4_921 (.A(\B_DOUT_TEMPR87[21] ), .B(\B_DOUT_TEMPR88[21] ), 
        .C(\B_DOUT_TEMPR89[21] ), .D(\B_DOUT_TEMPR90[21] ), .Y(
        OR4_921_Y));
    OR4 OR4_1225 (.A(\B_DOUT_TEMPR28[20] ), .B(\B_DOUT_TEMPR29[20] ), 
        .C(\B_DOUT_TEMPR30[20] ), .D(\B_DOUT_TEMPR31[20] ), .Y(
        OR4_1225_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%74%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R74C5 (
        .A_DOUT({nc16020, nc16021, nc16022, nc16023, nc16024, nc16025, 
        nc16026, nc16027, nc16028, nc16029, nc16030, nc16031, nc16032, 
        nc16033, nc16034, \A_DOUT_TEMPR74[29] , \A_DOUT_TEMPR74[28] , 
        \A_DOUT_TEMPR74[27] , \A_DOUT_TEMPR74[26] , 
        \A_DOUT_TEMPR74[25] }), .B_DOUT({nc16035, nc16036, nc16037, 
        nc16038, nc16039, nc16040, nc16041, nc16042, nc16043, nc16044, 
        nc16045, nc16046, nc16047, nc16048, nc16049, 
        \B_DOUT_TEMPR74[29] , \B_DOUT_TEMPR74[28] , 
        \B_DOUT_TEMPR74[27] , \B_DOUT_TEMPR74[26] , 
        \B_DOUT_TEMPR74[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[74][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1515 (.A(\A_DOUT_TEMPR79[0] ), .B(\A_DOUT_TEMPR80[0] ), .C(
        \A_DOUT_TEMPR81[0] ), .D(\A_DOUT_TEMPR82[0] ), .Y(OR4_1515_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%104%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R104C2 (
        .A_DOUT({nc16050, nc16051, nc16052, nc16053, nc16054, nc16055, 
        nc16056, nc16057, nc16058, nc16059, nc16060, nc16061, nc16062, 
        nc16063, nc16064, \A_DOUT_TEMPR104[14] , \A_DOUT_TEMPR104[13] , 
        \A_DOUT_TEMPR104[12] , \A_DOUT_TEMPR104[11] , 
        \A_DOUT_TEMPR104[10] }), .B_DOUT({nc16065, nc16066, nc16067, 
        nc16068, nc16069, nc16070, nc16071, nc16072, nc16073, nc16074, 
        nc16075, nc16076, nc16077, nc16078, nc16079, 
        \B_DOUT_TEMPR104[14] , \B_DOUT_TEMPR104[13] , 
        \B_DOUT_TEMPR104[12] , \B_DOUT_TEMPR104[11] , 
        \B_DOUT_TEMPR104[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[104][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_59 (.A(\A_DOUT_TEMPR72[24] ), .B(\A_DOUT_TEMPR73[24] ), .Y(
        OR2_59_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%93%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R93C6 (
        .A_DOUT({nc16080, nc16081, nc16082, nc16083, nc16084, nc16085, 
        nc16086, nc16087, nc16088, nc16089, nc16090, nc16091, nc16092, 
        nc16093, nc16094, \A_DOUT_TEMPR93[34] , \A_DOUT_TEMPR93[33] , 
        \A_DOUT_TEMPR93[32] , \A_DOUT_TEMPR93[31] , 
        \A_DOUT_TEMPR93[30] }), .B_DOUT({nc16095, nc16096, nc16097, 
        nc16098, nc16099, nc16100, nc16101, nc16102, nc16103, nc16104, 
        nc16105, nc16106, nc16107, nc16108, nc16109, 
        \B_DOUT_TEMPR93[34] , \B_DOUT_TEMPR93[33] , 
        \B_DOUT_TEMPR93[32] , \B_DOUT_TEMPR93[31] , 
        \B_DOUT_TEMPR93[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[93][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_302 (.A(\B_DOUT_TEMPR64[37] ), .B(\B_DOUT_TEMPR65[37] ), 
        .C(\B_DOUT_TEMPR66[37] ), .D(\B_DOUT_TEMPR67[37] ), .Y(
        OR4_302_Y));
    OR4 OR4_1784 (.A(OR4_540_Y), .B(OR4_852_Y), .C(OR4_474_Y), .D(
        OR4_876_Y), .Y(OR4_1784_Y));
    OR4 OR4_285 (.A(\B_DOUT_TEMPR79[10] ), .B(\B_DOUT_TEMPR80[10] ), 
        .C(\B_DOUT_TEMPR81[10] ), .D(\B_DOUT_TEMPR82[10] ), .Y(
        OR4_285_Y));
    OR4 OR4_2512 (.A(\A_DOUT_TEMPR79[23] ), .B(\A_DOUT_TEMPR80[23] ), 
        .C(\A_DOUT_TEMPR81[23] ), .D(\A_DOUT_TEMPR82[23] ), .Y(
        OR4_2512_Y));
    OR4 OR4_1481 (.A(\A_DOUT_TEMPR36[7] ), .B(\A_DOUT_TEMPR37[7] ), .C(
        \A_DOUT_TEMPR38[7] ), .D(\A_DOUT_TEMPR39[7] ), .Y(OR4_1481_Y));
    OR4 OR4_2623 (.A(\B_DOUT_TEMPR68[5] ), .B(\B_DOUT_TEMPR69[5] ), .C(
        \B_DOUT_TEMPR70[5] ), .D(\B_DOUT_TEMPR71[5] ), .Y(OR4_2623_Y));
    OR4 OR4_2404 (.A(OR4_2957_Y), .B(OR4_1239_Y), .C(OR4_878_Y), .D(
        OR4_1910_Y), .Y(OR4_2404_Y));
    OR4 OR4_1997 (.A(\B_DOUT_TEMPR107[6] ), .B(\B_DOUT_TEMPR108[6] ), 
        .C(\B_DOUT_TEMPR109[6] ), .D(\B_DOUT_TEMPR110[6] ), .Y(
        OR4_1997_Y));
    OR4 OR4_140 (.A(\A_DOUT_TEMPR83[0] ), .B(\A_DOUT_TEMPR84[0] ), .C(
        \A_DOUT_TEMPR85[0] ), .D(\A_DOUT_TEMPR86[0] ), .Y(OR4_140_Y));
    OR4 OR4_2781 (.A(\A_DOUT_TEMPR48[12] ), .B(\A_DOUT_TEMPR49[12] ), 
        .C(\A_DOUT_TEMPR50[12] ), .D(\A_DOUT_TEMPR51[12] ), .Y(
        OR4_2781_Y));
    OR4 OR4_2929 (.A(\B_DOUT_TEMPR0[3] ), .B(\B_DOUT_TEMPR1[3] ), .C(
        \B_DOUT_TEMPR2[3] ), .D(\B_DOUT_TEMPR3[3] ), .Y(OR4_2929_Y));
    OR4 OR4_686 (.A(\B_DOUT_TEMPR36[33] ), .B(\B_DOUT_TEMPR37[33] ), 
        .C(\B_DOUT_TEMPR38[33] ), .D(\B_DOUT_TEMPR39[33] ), .Y(
        OR4_686_Y));
    OR4 OR4_692 (.A(\A_DOUT_TEMPR60[23] ), .B(\A_DOUT_TEMPR61[23] ), 
        .C(\A_DOUT_TEMPR62[23] ), .D(\A_DOUT_TEMPR63[23] ), .Y(
        OR4_692_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%67%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R67C1 (
        .A_DOUT({nc16110, nc16111, nc16112, nc16113, nc16114, nc16115, 
        nc16116, nc16117, nc16118, nc16119, nc16120, nc16121, nc16122, 
        nc16123, nc16124, \A_DOUT_TEMPR67[9] , \A_DOUT_TEMPR67[8] , 
        \A_DOUT_TEMPR67[7] , \A_DOUT_TEMPR67[6] , \A_DOUT_TEMPR67[5] })
        , .B_DOUT({nc16125, nc16126, nc16127, nc16128, nc16129, 
        nc16130, nc16131, nc16132, nc16133, nc16134, nc16135, nc16136, 
        nc16137, nc16138, nc16139, \B_DOUT_TEMPR67[9] , 
        \B_DOUT_TEMPR67[8] , \B_DOUT_TEMPR67[7] , \B_DOUT_TEMPR67[6] , 
        \B_DOUT_TEMPR67[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[67][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_533 (.A(OR4_1943_Y), .B(OR4_1280_Y), .C(OR2_4_Y), .D(
        \B_DOUT_TEMPR74[0] ), .Y(OR4_533_Y));
    OR4 OR4_1049 (.A(\A_DOUT_TEMPR52[31] ), .B(\A_DOUT_TEMPR53[31] ), 
        .C(\A_DOUT_TEMPR54[31] ), .D(\A_DOUT_TEMPR55[31] ), .Y(
        OR4_1049_Y));
    OR4 OR4_2132 (.A(\B_DOUT_TEMPR75[17] ), .B(\B_DOUT_TEMPR76[17] ), 
        .C(\B_DOUT_TEMPR77[17] ), .D(\B_DOUT_TEMPR78[17] ), .Y(
        OR4_2132_Y));
    OR4 OR4_1805 (.A(\A_DOUT_TEMPR56[15] ), .B(\A_DOUT_TEMPR57[15] ), 
        .C(\A_DOUT_TEMPR58[15] ), .D(\A_DOUT_TEMPR59[15] ), .Y(
        OR4_1805_Y));
    OR4 OR4_2555 (.A(\B_DOUT_TEMPR64[38] ), .B(\B_DOUT_TEMPR65[38] ), 
        .C(\B_DOUT_TEMPR66[38] ), .D(\B_DOUT_TEMPR67[38] ), .Y(
        OR4_2555_Y));
    OR4 \OR4_B_DOUT[17]  (.A(OR4_2293_Y), .B(OR4_236_Y), .C(OR4_350_Y), 
        .D(OR4_231_Y), .Y(B_DOUT[17]));
    OR4 OR4_1549 (.A(\A_DOUT_TEMPR83[33] ), .B(\A_DOUT_TEMPR84[33] ), 
        .C(\A_DOUT_TEMPR85[33] ), .D(\A_DOUT_TEMPR86[33] ), .Y(
        OR4_1549_Y));
    OR4 OR4_2493 (.A(\A_DOUT_TEMPR20[31] ), .B(\A_DOUT_TEMPR21[31] ), 
        .C(\A_DOUT_TEMPR22[31] ), .D(\A_DOUT_TEMPR23[31] ), .Y(
        OR4_2493_Y));
    OR4 OR4_1132 (.A(\A_DOUT_TEMPR68[0] ), .B(\A_DOUT_TEMPR69[0] ), .C(
        \A_DOUT_TEMPR70[0] ), .D(\A_DOUT_TEMPR71[0] ), .Y(OR4_1132_Y));
    OR4 OR4_2074 (.A(\B_DOUT_TEMPR48[20] ), .B(\B_DOUT_TEMPR49[20] ), 
        .C(\B_DOUT_TEMPR50[20] ), .D(\B_DOUT_TEMPR51[20] ), .Y(
        OR4_2074_Y));
    OR4 OR4_1918 (.A(\A_DOUT_TEMPR12[5] ), .B(\A_DOUT_TEMPR13[5] ), .C(
        \A_DOUT_TEMPR14[5] ), .D(\A_DOUT_TEMPR15[5] ), .Y(OR4_1918_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%100%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R100C7 (
        .A_DOUT({nc16140, nc16141, nc16142, nc16143, nc16144, nc16145, 
        nc16146, nc16147, nc16148, nc16149, nc16150, nc16151, nc16152, 
        nc16153, nc16154, \A_DOUT_TEMPR100[39] , \A_DOUT_TEMPR100[38] , 
        \A_DOUT_TEMPR100[37] , \A_DOUT_TEMPR100[36] , 
        \A_DOUT_TEMPR100[35] }), .B_DOUT({nc16155, nc16156, nc16157, 
        nc16158, nc16159, nc16160, nc16161, nc16162, nc16163, nc16164, 
        nc16165, nc16166, nc16167, nc16168, nc16169, 
        \B_DOUT_TEMPR100[39] , \B_DOUT_TEMPR100[38] , 
        \B_DOUT_TEMPR100[37] , \B_DOUT_TEMPR100[36] , 
        \B_DOUT_TEMPR100[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[100][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_648 (.A(\B_DOUT_TEMPR16[14] ), .B(\B_DOUT_TEMPR17[14] ), 
        .C(\B_DOUT_TEMPR18[14] ), .D(\B_DOUT_TEMPR19[14] ), .Y(
        OR4_648_Y));
    OR4 OR4_2076 (.A(\B_DOUT_TEMPR111[17] ), .B(\B_DOUT_TEMPR112[17] ), 
        .C(\B_DOUT_TEMPR113[17] ), .D(\B_DOUT_TEMPR114[17] ), .Y(
        OR4_2076_Y));
    OR4 OR4_505 (.A(\B_DOUT_TEMPR99[27] ), .B(\B_DOUT_TEMPR100[27] ), 
        .C(\B_DOUT_TEMPR101[27] ), .D(\B_DOUT_TEMPR102[27] ), .Y(
        OR4_505_Y));
    OR4 OR4_924 (.A(OR4_530_Y), .B(OR4_1707_Y), .C(OR4_2796_Y), .D(
        OR4_1710_Y), .Y(OR4_924_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%31%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R31C0 (
        .A_DOUT({nc16170, nc16171, nc16172, nc16173, nc16174, nc16175, 
        nc16176, nc16177, nc16178, nc16179, nc16180, nc16181, nc16182, 
        nc16183, nc16184, \A_DOUT_TEMPR31[4] , \A_DOUT_TEMPR31[3] , 
        \A_DOUT_TEMPR31[2] , \A_DOUT_TEMPR31[1] , \A_DOUT_TEMPR31[0] })
        , .B_DOUT({nc16185, nc16186, nc16187, nc16188, nc16189, 
        nc16190, nc16191, nc16192, nc16193, nc16194, nc16195, nc16196, 
        nc16197, nc16198, nc16199, \B_DOUT_TEMPR31[4] , 
        \B_DOUT_TEMPR31[3] , \B_DOUT_TEMPR31[2] , \B_DOUT_TEMPR31[1] , 
        \B_DOUT_TEMPR31[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[22]  (.A(OR4_2300_Y), .B(OR4_901_Y), .C(OR4_1830_Y)
        , .D(OR4_1501_Y), .Y(A_DOUT[22]));
    OR4 OR4_1984 (.A(OR4_1874_Y), .B(OR4_492_Y), .C(OR4_1204_Y), .D(
        OR4_1472_Y), .Y(OR4_1984_Y));
    OR4 OR4_2724 (.A(\A_DOUT_TEMPR40[37] ), .B(\A_DOUT_TEMPR41[37] ), 
        .C(\A_DOUT_TEMPR42[37] ), .D(\A_DOUT_TEMPR43[37] ), .Y(
        OR4_2724_Y));
    OR4 OR4_1890 (.A(OR4_1628_Y), .B(OR4_2030_Y), .C(OR4_2794_Y), .D(
        OR4_549_Y), .Y(OR4_1890_Y));
    OR2 OR2_36 (.A(\B_DOUT_TEMPR72[5] ), .B(\B_DOUT_TEMPR73[5] ), .Y(
        OR2_36_Y));
    OR4 OR4_1342 (.A(OR4_41_Y), .B(OR4_2312_Y), .C(OR4_761_Y), .D(
        OR4_2313_Y), .Y(OR4_1342_Y));
    OR4 OR4_2421 (.A(\B_DOUT_TEMPR44[18] ), .B(\B_DOUT_TEMPR45[18] ), 
        .C(\B_DOUT_TEMPR46[18] ), .D(\B_DOUT_TEMPR47[18] ), .Y(
        OR4_2421_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%102%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R102C4 (
        .A_DOUT({nc16200, nc16201, nc16202, nc16203, nc16204, nc16205, 
        nc16206, nc16207, nc16208, nc16209, nc16210, nc16211, nc16212, 
        nc16213, nc16214, \A_DOUT_TEMPR102[24] , \A_DOUT_TEMPR102[23] , 
        \A_DOUT_TEMPR102[22] , \A_DOUT_TEMPR102[21] , 
        \A_DOUT_TEMPR102[20] }), .B_DOUT({nc16215, nc16216, nc16217, 
        nc16218, nc16219, nc16220, nc16221, nc16222, nc16223, nc16224, 
        nc16225, nc16226, nc16227, nc16228, nc16229, 
        \B_DOUT_TEMPR102[24] , \B_DOUT_TEMPR102[23] , 
        \B_DOUT_TEMPR102[22] , \B_DOUT_TEMPR102[21] , 
        \B_DOUT_TEMPR102[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[102][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1986 (.A(OR4_1122_Y), .B(OR4_2799_Y), .C(OR4_2137_Y), .D(
        OR4_1466_Y), .Y(OR4_1986_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%94%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R94C4 (
        .A_DOUT({nc16230, nc16231, nc16232, nc16233, nc16234, nc16235, 
        nc16236, nc16237, nc16238, nc16239, nc16240, nc16241, nc16242, 
        nc16243, nc16244, \A_DOUT_TEMPR94[24] , \A_DOUT_TEMPR94[23] , 
        \A_DOUT_TEMPR94[22] , \A_DOUT_TEMPR94[21] , 
        \A_DOUT_TEMPR94[20] }), .B_DOUT({nc16245, nc16246, nc16247, 
        nc16248, nc16249, nc16250, nc16251, nc16252, nc16253, nc16254, 
        nc16255, nc16256, nc16257, nc16258, nc16259, 
        \B_DOUT_TEMPR94[24] , \B_DOUT_TEMPR94[23] , 
        \B_DOUT_TEMPR94[22] , \B_DOUT_TEMPR94[21] , 
        \B_DOUT_TEMPR94[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[94][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_941 (.A(\B_DOUT_TEMPR95[31] ), .B(\B_DOUT_TEMPR96[31] ), 
        .C(\B_DOUT_TEMPR97[31] ), .D(\B_DOUT_TEMPR98[31] ), .Y(
        OR4_941_Y));
    OR4 OR4_1771 (.A(\B_DOUT_TEMPR16[38] ), .B(\B_DOUT_TEMPR17[38] ), 
        .C(\B_DOUT_TEMPR18[38] ), .D(\B_DOUT_TEMPR19[38] ), .Y(
        OR4_1771_Y));
    OR4 OR4_1054 (.A(OR4_451_Y), .B(OR4_1766_Y), .C(OR4_1417_Y), .D(
        OR4_2464_Y), .Y(OR4_1054_Y));
    OR4 OR4_2373 (.A(\A_DOUT_TEMPR60[6] ), .B(\A_DOUT_TEMPR61[6] ), .C(
        \A_DOUT_TEMPR62[6] ), .D(\A_DOUT_TEMPR63[6] ), .Y(OR4_2373_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%5%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R5C0 (
        .A_DOUT({nc16260, nc16261, nc16262, nc16263, nc16264, nc16265, 
        nc16266, nc16267, nc16268, nc16269, nc16270, nc16271, nc16272, 
        nc16273, nc16274, \A_DOUT_TEMPR5[4] , \A_DOUT_TEMPR5[3] , 
        \A_DOUT_TEMPR5[2] , \A_DOUT_TEMPR5[1] , \A_DOUT_TEMPR5[0] }), 
        .B_DOUT({nc16275, nc16276, nc16277, nc16278, nc16279, nc16280, 
        nc16281, nc16282, nc16283, nc16284, nc16285, nc16286, nc16287, 
        nc16288, nc16289, \B_DOUT_TEMPR5[4] , \B_DOUT_TEMPR5[3] , 
        \B_DOUT_TEMPR5[2] , \B_DOUT_TEMPR5[1] , \B_DOUT_TEMPR5[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[5][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[1] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[1] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%89%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R89C3 (
        .A_DOUT({nc16290, nc16291, nc16292, nc16293, nc16294, nc16295, 
        nc16296, nc16297, nc16298, nc16299, nc16300, nc16301, nc16302, 
        nc16303, nc16304, \A_DOUT_TEMPR89[19] , \A_DOUT_TEMPR89[18] , 
        \A_DOUT_TEMPR89[17] , \A_DOUT_TEMPR89[16] , 
        \A_DOUT_TEMPR89[15] }), .B_DOUT({nc16305, nc16306, nc16307, 
        nc16308, nc16309, nc16310, nc16311, nc16312, nc16313, nc16314, 
        nc16315, nc16316, nc16317, nc16318, nc16319, 
        \B_DOUT_TEMPR89[19] , \B_DOUT_TEMPR89[18] , 
        \B_DOUT_TEMPR89[17] , \B_DOUT_TEMPR89[16] , 
        \B_DOUT_TEMPR89[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[89][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1894 (.A(OR4_2436_Y), .B(OR4_310_Y), .C(OR4_3024_Y), .D(
        OR4_1459_Y), .Y(OR4_1894_Y));
    OR4 OR4_184 (.A(OR4_1964_Y), .B(OR4_777_Y), .C(OR4_2239_Y), .D(
        OR4_779_Y), .Y(OR4_184_Y));
    OR4 OR4_1056 (.A(\A_DOUT_TEMPR16[12] ), .B(\A_DOUT_TEMPR17[12] ), 
        .C(\A_DOUT_TEMPR18[12] ), .D(\A_DOUT_TEMPR19[12] ), .Y(
        OR4_1056_Y));
    OR4 OR4_384 (.A(OR4_1827_Y), .B(OR4_1166_Y), .C(OR4_714_Y), .D(
        OR4_2383_Y), .Y(OR4_384_Y));
    OR4 OR4_2483 (.A(\B_DOUT_TEMPR60[35] ), .B(\B_DOUT_TEMPR61[35] ), 
        .C(\B_DOUT_TEMPR62[35] ), .D(\B_DOUT_TEMPR63[35] ), .Y(
        OR4_2483_Y));
    OR4 OR4_1564 (.A(\B_DOUT_TEMPR83[14] ), .B(\B_DOUT_TEMPR84[14] ), 
        .C(\B_DOUT_TEMPR85[14] ), .D(\B_DOUT_TEMPR86[14] ), .Y(
        OR4_1564_Y));
    OR4 OR4_2010 (.A(\A_DOUT_TEMPR36[37] ), .B(\A_DOUT_TEMPR37[37] ), 
        .C(\A_DOUT_TEMPR38[37] ), .D(\A_DOUT_TEMPR39[37] ), .Y(
        OR4_2010_Y));
    OR4 OR4_2958 (.A(\A_DOUT_TEMPR24[4] ), .B(\A_DOUT_TEMPR25[4] ), .C(
        \A_DOUT_TEMPR26[4] ), .D(\A_DOUT_TEMPR27[4] ), .Y(OR4_2958_Y));
    OR4 OR4_1626 (.A(OR4_1787_Y), .B(OR4_1136_Y), .C(OR4_17_Y), .D(
        OR4_2364_Y), .Y(OR4_1626_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%78%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R78C4 (
        .A_DOUT({nc16320, nc16321, nc16322, nc16323, nc16324, nc16325, 
        nc16326, nc16327, nc16328, nc16329, nc16330, nc16331, nc16332, 
        nc16333, nc16334, \A_DOUT_TEMPR78[24] , \A_DOUT_TEMPR78[23] , 
        \A_DOUT_TEMPR78[22] , \A_DOUT_TEMPR78[21] , 
        \A_DOUT_TEMPR78[20] }), .B_DOUT({nc16335, nc16336, nc16337, 
        nc16338, nc16339, nc16340, nc16341, nc16342, nc16343, nc16344, 
        nc16345, nc16346, nc16347, nc16348, nc16349, 
        \B_DOUT_TEMPR78[24] , \B_DOUT_TEMPR78[23] , 
        \B_DOUT_TEMPR78[22] , \B_DOUT_TEMPR78[21] , 
        \B_DOUT_TEMPR78[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[78][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%43%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R43C4 (
        .A_DOUT({nc16350, nc16351, nc16352, nc16353, nc16354, nc16355, 
        nc16356, nc16357, nc16358, nc16359, nc16360, nc16361, nc16362, 
        nc16363, nc16364, \A_DOUT_TEMPR43[24] , \A_DOUT_TEMPR43[23] , 
        \A_DOUT_TEMPR43[22] , \A_DOUT_TEMPR43[21] , 
        \A_DOUT_TEMPR43[20] }), .B_DOUT({nc16365, nc16366, nc16367, 
        nc16368, nc16369, nc16370, nc16371, nc16372, nc16373, nc16374, 
        nc16375, nc16376, nc16377, nc16378, nc16379, 
        \B_DOUT_TEMPR43[24] , \B_DOUT_TEMPR43[23] , 
        \B_DOUT_TEMPR43[22] , \B_DOUT_TEMPR43[21] , 
        \B_DOUT_TEMPR43[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[43][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1120 (.A(\B_DOUT_TEMPR91[5] ), .B(\B_DOUT_TEMPR92[5] ), .C(
        \B_DOUT_TEMPR93[5] ), .D(\B_DOUT_TEMPR94[5] ), .Y(OR4_1120_Y));
    OR4 OR4_2204 (.A(\B_DOUT_TEMPR36[1] ), .B(\B_DOUT_TEMPR37[1] ), .C(
        \B_DOUT_TEMPR38[1] ), .D(\B_DOUT_TEMPR39[1] ), .Y(OR4_2204_Y));
    OR4 OR4_1117 (.A(\A_DOUT_TEMPR99[19] ), .B(\A_DOUT_TEMPR100[19] ), 
        .C(\A_DOUT_TEMPR101[19] ), .D(\A_DOUT_TEMPR102[19] ), .Y(
        OR4_1117_Y));
    OR4 OR4_463 (.A(\A_DOUT_TEMPR12[37] ), .B(\A_DOUT_TEMPR13[37] ), 
        .C(\A_DOUT_TEMPR14[37] ), .D(\A_DOUT_TEMPR15[37] ), .Y(
        OR4_463_Y));
    OR4 OR4_1614 (.A(\A_DOUT_TEMPR24[1] ), .B(\A_DOUT_TEMPR25[1] ), .C(
        \A_DOUT_TEMPR26[1] ), .D(\A_DOUT_TEMPR27[1] ), .Y(OR4_1614_Y));
    OR4 OR4_1353 (.A(\A_DOUT_TEMPR48[2] ), .B(\A_DOUT_TEMPR49[2] ), .C(
        \A_DOUT_TEMPR50[2] ), .D(\A_DOUT_TEMPR51[2] ), .Y(OR4_1353_Y));
    OR4 OR4_352 (.A(\A_DOUT_TEMPR8[10] ), .B(\A_DOUT_TEMPR9[10] ), .C(
        \A_DOUT_TEMPR10[10] ), .D(\A_DOUT_TEMPR11[10] ), .Y(OR4_352_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%87%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R87C3 (
        .A_DOUT({nc16380, nc16381, nc16382, nc16383, nc16384, nc16385, 
        nc16386, nc16387, nc16388, nc16389, nc16390, nc16391, nc16392, 
        nc16393, nc16394, \A_DOUT_TEMPR87[19] , \A_DOUT_TEMPR87[18] , 
        \A_DOUT_TEMPR87[17] , \A_DOUT_TEMPR87[16] , 
        \A_DOUT_TEMPR87[15] }), .B_DOUT({nc16395, nc16396, nc16397, 
        nc16398, nc16399, nc16400, nc16401, nc16402, nc16403, nc16404, 
        nc16405, nc16406, nc16407, nc16408, nc16409, 
        \B_DOUT_TEMPR87[19] , \B_DOUT_TEMPR87[18] , 
        \B_DOUT_TEMPR87[17] , \B_DOUT_TEMPR87[16] , 
        \B_DOUT_TEMPR87[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[87][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1545 (.A(OR4_2080_Y), .B(OR4_2961_Y), .C(OR4_1391_Y), .D(
        OR4_2963_Y), .Y(OR4_1545_Y));
    OR4 OR4_2924 (.A(\B_DOUT_TEMPR8[29] ), .B(\B_DOUT_TEMPR9[29] ), .C(
        \B_DOUT_TEMPR10[29] ), .D(\B_DOUT_TEMPR11[29] ), .Y(OR4_2924_Y)
        );
    CFG3 #( .INIT(8'h8) )  CFG3_19 (.A(B_ADDR[16]), .B(B_ADDR[15]), .C(
        B_ADDR[14]), .Y(CFG3_19_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%7%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R7C0 (
        .A_DOUT({nc16410, nc16411, nc16412, nc16413, nc16414, nc16415, 
        nc16416, nc16417, nc16418, nc16419, nc16420, nc16421, nc16422, 
        nc16423, nc16424, \A_DOUT_TEMPR7[4] , \A_DOUT_TEMPR7[3] , 
        \A_DOUT_TEMPR7[2] , \A_DOUT_TEMPR7[1] , \A_DOUT_TEMPR7[0] }), 
        .B_DOUT({nc16425, nc16426, nc16427, nc16428, nc16429, nc16430, 
        nc16431, nc16432, nc16433, nc16434, nc16435, nc16436, nc16437, 
        nc16438, nc16439, \B_DOUT_TEMPR7[4] , \B_DOUT_TEMPR7[3] , 
        \B_DOUT_TEMPR7[2] , \B_DOUT_TEMPR7[1] , \B_DOUT_TEMPR7[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[7][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[1] , A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[1] , B_ADDR[13], B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%19%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R19C6 (
        .A_DOUT({nc16440, nc16441, nc16442, nc16443, nc16444, nc16445, 
        nc16446, nc16447, nc16448, nc16449, nc16450, nc16451, nc16452, 
        nc16453, nc16454, \A_DOUT_TEMPR19[34] , \A_DOUT_TEMPR19[33] , 
        \A_DOUT_TEMPR19[32] , \A_DOUT_TEMPR19[31] , 
        \A_DOUT_TEMPR19[30] }), .B_DOUT({nc16455, nc16456, nc16457, 
        nc16458, nc16459, nc16460, nc16461, nc16462, nc16463, nc16464, 
        nc16465, nc16466, nc16467, nc16468, nc16469, 
        \B_DOUT_TEMPR19[34] , \B_DOUT_TEMPR19[33] , 
        \B_DOUT_TEMPR19[32] , \B_DOUT_TEMPR19[31] , 
        \B_DOUT_TEMPR19[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2003 (.A(\B_DOUT_TEMPR0[12] ), .B(\B_DOUT_TEMPR1[12] ), .C(
        \B_DOUT_TEMPR2[12] ), .D(\B_DOUT_TEMPR3[12] ), .Y(OR4_2003_Y));
    OR4 OR4_1261 (.A(\A_DOUT_TEMPR99[28] ), .B(\A_DOUT_TEMPR100[28] ), 
        .C(\A_DOUT_TEMPR101[28] ), .D(\A_DOUT_TEMPR102[28] ), .Y(
        OR4_1261_Y));
    OR4 OR4_2926 (.A(\B_DOUT_TEMPR103[32] ), .B(\B_DOUT_TEMPR104[32] ), 
        .C(\B_DOUT_TEMPR105[32] ), .D(\B_DOUT_TEMPR106[32] ), .Y(
        OR4_2926_Y));
    OR4 OR4_2601 (.A(\A_DOUT_TEMPR115[3] ), .B(\A_DOUT_TEMPR116[3] ), 
        .C(\A_DOUT_TEMPR117[3] ), .D(\A_DOUT_TEMPR118[3] ), .Y(
        OR4_2601_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%105%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R105C4 (
        .A_DOUT({nc16470, nc16471, nc16472, nc16473, nc16474, nc16475, 
        nc16476, nc16477, nc16478, nc16479, nc16480, nc16481, nc16482, 
        nc16483, nc16484, \A_DOUT_TEMPR105[24] , \A_DOUT_TEMPR105[23] , 
        \A_DOUT_TEMPR105[22] , \A_DOUT_TEMPR105[21] , 
        \A_DOUT_TEMPR105[20] }), .B_DOUT({nc16485, nc16486, nc16487, 
        nc16488, nc16489, nc16490, nc16491, nc16492, nc16493, nc16494, 
        nc16495, nc16496, nc16497, nc16498, nc16499, 
        \B_DOUT_TEMPR105[24] , \B_DOUT_TEMPR105[23] , 
        \B_DOUT_TEMPR105[22] , \B_DOUT_TEMPR105[21] , 
        \B_DOUT_TEMPR105[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[105][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[28]  (.A(CFG3_12_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[28] ));
    OR4 OR4_944 (.A(\A_DOUT_TEMPR28[16] ), .B(\A_DOUT_TEMPR29[16] ), 
        .C(\A_DOUT_TEMPR30[16] ), .D(\A_DOUT_TEMPR31[16] ), .Y(
        OR4_944_Y));
    OR4 OR4_1473 (.A(\B_DOUT_TEMPR107[24] ), .B(\B_DOUT_TEMPR108[24] ), 
        .C(\B_DOUT_TEMPR109[24] ), .D(\B_DOUT_TEMPR110[24] ), .Y(
        OR4_1473_Y));
    OR4 OR4_3009 (.A(\A_DOUT_TEMPR115[36] ), .B(\A_DOUT_TEMPR116[36] ), 
        .C(\A_DOUT_TEMPR117[36] ), .D(\A_DOUT_TEMPR118[36] ), .Y(
        OR4_3009_Y));
    OR4 OR4_2703 (.A(\B_DOUT_TEMPR103[38] ), .B(\B_DOUT_TEMPR104[38] ), 
        .C(\B_DOUT_TEMPR105[38] ), .D(\B_DOUT_TEMPR106[38] ), .Y(
        OR4_2703_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%57%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R57C4 (
        .A_DOUT({nc16500, nc16501, nc16502, nc16503, nc16504, nc16505, 
        nc16506, nc16507, nc16508, nc16509, nc16510, nc16511, nc16512, 
        nc16513, nc16514, \A_DOUT_TEMPR57[24] , \A_DOUT_TEMPR57[23] , 
        \A_DOUT_TEMPR57[22] , \A_DOUT_TEMPR57[21] , 
        \A_DOUT_TEMPR57[20] }), .B_DOUT({nc16515, nc16516, nc16517, 
        nc16518, nc16519, nc16520, nc16521, nc16522, nc16523, nc16524, 
        nc16525, nc16526, nc16527, nc16528, nc16529, 
        \B_DOUT_TEMPR57[24] , \B_DOUT_TEMPR57[23] , 
        \B_DOUT_TEMPR57[22] , \B_DOUT_TEMPR57[21] , 
        \B_DOUT_TEMPR57[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[57][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_72 (.A(\A_DOUT_TEMPR72[26] ), .B(\A_DOUT_TEMPR73[26] ), .Y(
        OR2_72_Y));
    OR4 OR4_2157 (.A(\A_DOUT_TEMPR48[7] ), .B(\A_DOUT_TEMPR49[7] ), .C(
        \A_DOUT_TEMPR50[7] ), .D(\A_DOUT_TEMPR51[7] ), .Y(OR4_2157_Y));
    OR4 OR4_2416 (.A(OR4_2802_Y), .B(OR4_1078_Y), .C(OR4_703_Y), .D(
        OR4_1741_Y), .Y(OR4_2416_Y));
    OR4 OR4_2654 (.A(OR4_2006_Y), .B(OR4_462_Y), .C(OR4_1066_Y), .D(
        OR4_868_Y), .Y(OR4_2654_Y));
    OR4 OR4_2105 (.A(\B_DOUT_TEMPR75[21] ), .B(\B_DOUT_TEMPR76[21] ), 
        .C(\B_DOUT_TEMPR77[21] ), .D(\B_DOUT_TEMPR78[21] ), .Y(
        OR4_2105_Y));
    OR4 OR4_410 (.A(\B_DOUT_TEMPR32[6] ), .B(\B_DOUT_TEMPR33[6] ), .C(
        \B_DOUT_TEMPR34[6] ), .D(\B_DOUT_TEMPR35[6] ), .Y(OR4_410_Y));
    OR4 OR4_378 (.A(\A_DOUT_TEMPR56[33] ), .B(\A_DOUT_TEMPR57[33] ), 
        .C(\A_DOUT_TEMPR58[33] ), .D(\A_DOUT_TEMPR59[33] ), .Y(
        OR4_378_Y));
    OR4 OR4_2239 (.A(\A_DOUT_TEMPR40[16] ), .B(\A_DOUT_TEMPR41[16] ), 
        .C(\A_DOUT_TEMPR42[16] ), .D(\A_DOUT_TEMPR43[16] ), .Y(
        OR4_2239_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%41%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R41C4 (
        .A_DOUT({nc16530, nc16531, nc16532, nc16533, nc16534, nc16535, 
        nc16536, nc16537, nc16538, nc16539, nc16540, nc16541, nc16542, 
        nc16543, nc16544, \A_DOUT_TEMPR41[24] , \A_DOUT_TEMPR41[23] , 
        \A_DOUT_TEMPR41[22] , \A_DOUT_TEMPR41[21] , 
        \A_DOUT_TEMPR41[20] }), .B_DOUT({nc16545, nc16546, nc16547, 
        nc16548, nc16549, nc16550, nc16551, nc16552, nc16553, nc16554, 
        nc16555, nc16556, nc16557, nc16558, nc16559, 
        \B_DOUT_TEMPR41[24] , \B_DOUT_TEMPR41[23] , 
        \B_DOUT_TEMPR41[22] , \B_DOUT_TEMPR41[21] , 
        \B_DOUT_TEMPR41[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[41][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_775 (.A(\A_DOUT_TEMPR20[19] ), .B(\A_DOUT_TEMPR21[19] ), 
        .C(\A_DOUT_TEMPR22[19] ), .D(\A_DOUT_TEMPR23[19] ), .Y(
        OR4_775_Y));
    OR4 OR4_555 (.A(\A_DOUT_TEMPR16[25] ), .B(\A_DOUT_TEMPR17[25] ), 
        .C(\A_DOUT_TEMPR18[25] ), .D(\A_DOUT_TEMPR19[25] ), .Y(
        OR4_555_Y));
    OR4 OR4_1948 (.A(\B_DOUT_TEMPR24[39] ), .B(\B_DOUT_TEMPR25[39] ), 
        .C(\B_DOUT_TEMPR26[39] ), .D(\B_DOUT_TEMPR27[39] ), .Y(
        OR4_1948_Y));
    OR4 OR4_2296 (.A(OR4_2453_Y), .B(OR4_1631_Y), .C(OR4_618_Y), .D(
        OR4_951_Y), .Y(OR4_2296_Y));
    OR4 OR4_1239 (.A(\A_DOUT_TEMPR91[5] ), .B(\A_DOUT_TEMPR92[5] ), .C(
        \A_DOUT_TEMPR93[5] ), .D(\A_DOUT_TEMPR94[5] ), .Y(OR4_1239_Y));
    OR4 OR4_886 (.A(\A_DOUT_TEMPR75[24] ), .B(\A_DOUT_TEMPR76[24] ), 
        .C(\A_DOUT_TEMPR77[24] ), .D(\A_DOUT_TEMPR78[24] ), .Y(
        OR4_886_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%53%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R53C6 (
        .A_DOUT({nc16560, nc16561, nc16562, nc16563, nc16564, nc16565, 
        nc16566, nc16567, nc16568, nc16569, nc16570, nc16571, nc16572, 
        nc16573, nc16574, \A_DOUT_TEMPR53[34] , \A_DOUT_TEMPR53[33] , 
        \A_DOUT_TEMPR53[32] , \A_DOUT_TEMPR53[31] , 
        \A_DOUT_TEMPR53[30] }), .B_DOUT({nc16575, nc16576, nc16577, 
        nc16578, nc16579, nc16580, nc16581, nc16582, nc16583, nc16584, 
        nc16585, nc16586, nc16587, nc16588, nc16589, 
        \B_DOUT_TEMPR53[34] , \B_DOUT_TEMPR53[33] , 
        \B_DOUT_TEMPR53[32] , \B_DOUT_TEMPR53[31] , 
        \B_DOUT_TEMPR53[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[53][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%74%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R74C7 (
        .A_DOUT({nc16590, nc16591, nc16592, nc16593, nc16594, nc16595, 
        nc16596, nc16597, nc16598, nc16599, nc16600, nc16601, nc16602, 
        nc16603, nc16604, \A_DOUT_TEMPR74[39] , \A_DOUT_TEMPR74[38] , 
        \A_DOUT_TEMPR74[37] , \A_DOUT_TEMPR74[36] , 
        \A_DOUT_TEMPR74[35] }), .B_DOUT({nc16605, nc16606, nc16607, 
        nc16608, nc16609, nc16610, nc16611, nc16612, nc16613, nc16614, 
        nc16615, nc16616, nc16617, nc16618, nc16619, 
        \B_DOUT_TEMPR74[39] , \B_DOUT_TEMPR74[38] , 
        \B_DOUT_TEMPR74[37] , \B_DOUT_TEMPR74[36] , 
        \B_DOUT_TEMPR74[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[74][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2715 (.A(\B_DOUT_TEMPR115[36] ), .B(\B_DOUT_TEMPR116[36] ), 
        .C(\B_DOUT_TEMPR117[36] ), .D(\B_DOUT_TEMPR118[36] ), .Y(
        OR4_2715_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%17%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R17C1 (
        .A_DOUT({nc16620, nc16621, nc16622, nc16623, nc16624, nc16625, 
        nc16626, nc16627, nc16628, nc16629, nc16630, nc16631, nc16632, 
        nc16633, nc16634, \A_DOUT_TEMPR17[9] , \A_DOUT_TEMPR17[8] , 
        \A_DOUT_TEMPR17[7] , \A_DOUT_TEMPR17[6] , \A_DOUT_TEMPR17[5] })
        , .B_DOUT({nc16635, nc16636, nc16637, nc16638, nc16639, 
        nc16640, nc16641, nc16642, nc16643, nc16644, nc16645, nc16646, 
        nc16647, nc16648, nc16649, \B_DOUT_TEMPR17[9] , 
        \B_DOUT_TEMPR17[8] , \B_DOUT_TEMPR17[7] , \B_DOUT_TEMPR17[6] , 
        \B_DOUT_TEMPR17[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2761 (.A(\A_DOUT_TEMPR36[10] ), .B(\A_DOUT_TEMPR37[10] ), 
        .C(\A_DOUT_TEMPR38[10] ), .D(\A_DOUT_TEMPR39[10] ), .Y(
        OR4_2761_Y));
    OR4 OR4_2001 (.A(\B_DOUT_TEMPR95[33] ), .B(\B_DOUT_TEMPR96[33] ), 
        .C(\B_DOUT_TEMPR97[33] ), .D(\B_DOUT_TEMPR98[33] ), .Y(
        OR4_2001_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_7 (.A(VCC), .B(A_ADDR[18]), .C(
        A_ADDR[17]), .Y(CFG3_7_Y));
    OR4 OR4_380 (.A(\B_DOUT_TEMPR68[29] ), .B(\B_DOUT_TEMPR69[29] ), 
        .C(\B_DOUT_TEMPR70[29] ), .D(\B_DOUT_TEMPR71[29] ), .Y(
        OR4_380_Y));
    OR4 OR4_1608 (.A(\A_DOUT_TEMPR12[24] ), .B(\A_DOUT_TEMPR13[24] ), 
        .C(\A_DOUT_TEMPR14[24] ), .D(\A_DOUT_TEMPR15[24] ), .Y(
        OR4_1608_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%41%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R41C3 (
        .A_DOUT({nc16650, nc16651, nc16652, nc16653, nc16654, nc16655, 
        nc16656, nc16657, nc16658, nc16659, nc16660, nc16661, nc16662, 
        nc16663, nc16664, \A_DOUT_TEMPR41[19] , \A_DOUT_TEMPR41[18] , 
        \A_DOUT_TEMPR41[17] , \A_DOUT_TEMPR41[16] , 
        \A_DOUT_TEMPR41[15] }), .B_DOUT({nc16665, nc16666, nc16667, 
        nc16668, nc16669, nc16670, nc16671, nc16672, nc16673, nc16674, 
        nc16675, nc16676, nc16677, nc16678, nc16679, 
        \B_DOUT_TEMPR41[19] , \B_DOUT_TEMPR41[18] , 
        \B_DOUT_TEMPR41[17] , \B_DOUT_TEMPR41[16] , 
        \B_DOUT_TEMPR41[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[41][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[1]  (.A(OR4_1532_Y), .B(OR4_1853_Y), .C(OR4_2716_Y)
        , .D(OR4_2773_Y), .Y(B_DOUT[1]));
    OR4 OR4_1923 (.A(\B_DOUT_TEMPR40[14] ), .B(\B_DOUT_TEMPR41[14] ), 
        .C(\B_DOUT_TEMPR42[14] ), .D(\B_DOUT_TEMPR43[14] ), .Y(
        OR4_1923_Y));
    OR4 OR4_978 (.A(\A_DOUT_TEMPR95[4] ), .B(\A_DOUT_TEMPR96[4] ), .C(
        \A_DOUT_TEMPR97[4] ), .D(\A_DOUT_TEMPR98[4] ), .Y(OR4_978_Y));
    OR4 OR4_2286 (.A(\B_DOUT_TEMPR60[18] ), .B(\B_DOUT_TEMPR61[18] ), 
        .C(\B_DOUT_TEMPR62[18] ), .D(\B_DOUT_TEMPR63[18] ), .Y(
        OR4_2286_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%61%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R61C0 (
        .A_DOUT({nc16680, nc16681, nc16682, nc16683, nc16684, nc16685, 
        nc16686, nc16687, nc16688, nc16689, nc16690, nc16691, nc16692, 
        nc16693, nc16694, \A_DOUT_TEMPR61[4] , \A_DOUT_TEMPR61[3] , 
        \A_DOUT_TEMPR61[2] , \A_DOUT_TEMPR61[1] , \A_DOUT_TEMPR61[0] })
        , .B_DOUT({nc16695, nc16696, nc16697, nc16698, nc16699, 
        nc16700, nc16701, nc16702, nc16703, nc16704, nc16705, nc16706, 
        nc16707, nc16708, nc16709, \B_DOUT_TEMPR61[4] , 
        \B_DOUT_TEMPR61[3] , \B_DOUT_TEMPR61[2] , \B_DOUT_TEMPR61[1] , 
        \B_DOUT_TEMPR61[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[61][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_429 (.A(OR4_2031_Y), .B(OR4_2019_Y), .C(OR4_2659_Y), .D(
        OR4_1831_Y), .Y(OR4_429_Y));
    OR4 OR4_1395 (.A(\A_DOUT_TEMPR0[11] ), .B(\A_DOUT_TEMPR1[11] ), .C(
        \A_DOUT_TEMPR2[11] ), .D(\A_DOUT_TEMPR3[11] ), .Y(OR4_1395_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%86%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R86C5 (
        .A_DOUT({nc16710, nc16711, nc16712, nc16713, nc16714, nc16715, 
        nc16716, nc16717, nc16718, nc16719, nc16720, nc16721, nc16722, 
        nc16723, nc16724, \A_DOUT_TEMPR86[29] , \A_DOUT_TEMPR86[28] , 
        \A_DOUT_TEMPR86[27] , \A_DOUT_TEMPR86[26] , 
        \A_DOUT_TEMPR86[25] }), .B_DOUT({nc16725, nc16726, nc16727, 
        nc16728, nc16729, nc16730, nc16731, nc16732, nc16733, nc16734, 
        nc16735, nc16736, nc16737, nc16738, nc16739, 
        \B_DOUT_TEMPR86[29] , \B_DOUT_TEMPR86[28] , 
        \B_DOUT_TEMPR86[27] , \B_DOUT_TEMPR86[26] , 
        \B_DOUT_TEMPR86[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[86][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%89%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R89C5 (
        .A_DOUT({nc16740, nc16741, nc16742, nc16743, nc16744, nc16745, 
        nc16746, nc16747, nc16748, nc16749, nc16750, nc16751, nc16752, 
        nc16753, nc16754, \A_DOUT_TEMPR89[29] , \A_DOUT_TEMPR89[28] , 
        \A_DOUT_TEMPR89[27] , \A_DOUT_TEMPR89[26] , 
        \A_DOUT_TEMPR89[25] }), .B_DOUT({nc16755, nc16756, nc16757, 
        nc16758, nc16759, nc16760, nc16761, nc16762, nc16763, nc16764, 
        nc16765, nc16766, nc16767, nc16768, nc16769, 
        \B_DOUT_TEMPR89[29] , \B_DOUT_TEMPR89[28] , 
        \B_DOUT_TEMPR89[27] , \B_DOUT_TEMPR89[26] , 
        \B_DOUT_TEMPR89[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[89][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_119 (.A(\B_DOUT_TEMPR24[3] ), .B(\B_DOUT_TEMPR25[3] ), .C(
        \B_DOUT_TEMPR26[3] ), .D(\B_DOUT_TEMPR27[3] ), .Y(OR4_119_Y));
    OR4 OR4_308 (.A(\B_DOUT_TEMPR91[35] ), .B(\B_DOUT_TEMPR92[35] ), 
        .C(\B_DOUT_TEMPR93[35] ), .D(\B_DOUT_TEMPR94[35] ), .Y(
        OR4_308_Y));
    OR4 OR4_1147 (.A(\A_DOUT_TEMPR24[26] ), .B(\A_DOUT_TEMPR25[26] ), 
        .C(\A_DOUT_TEMPR26[26] ), .D(\A_DOUT_TEMPR27[26] ), .Y(
        OR4_1147_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%37%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R37C4 (
        .A_DOUT({nc16770, nc16771, nc16772, nc16773, nc16774, nc16775, 
        nc16776, nc16777, nc16778, nc16779, nc16780, nc16781, nc16782, 
        nc16783, nc16784, \A_DOUT_TEMPR37[24] , \A_DOUT_TEMPR37[23] , 
        \A_DOUT_TEMPR37[22] , \A_DOUT_TEMPR37[21] , 
        \A_DOUT_TEMPR37[20] }), .B_DOUT({nc16785, nc16786, nc16787, 
        nc16788, nc16789, nc16790, nc16791, nc16792, nc16793, nc16794, 
        nc16795, nc16796, nc16797, nc16798, nc16799, 
        \B_DOUT_TEMPR37[24] , \B_DOUT_TEMPR37[23] , 
        \B_DOUT_TEMPR37[22] , \B_DOUT_TEMPR37[21] , 
        \B_DOUT_TEMPR37[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[37][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%92%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R92C7 (
        .A_DOUT({nc16800, nc16801, nc16802, nc16803, nc16804, nc16805, 
        nc16806, nc16807, nc16808, nc16809, nc16810, nc16811, nc16812, 
        nc16813, nc16814, \A_DOUT_TEMPR92[39] , \A_DOUT_TEMPR92[38] , 
        \A_DOUT_TEMPR92[37] , \A_DOUT_TEMPR92[36] , 
        \A_DOUT_TEMPR92[35] }), .B_DOUT({nc16815, nc16816, nc16817, 
        nc16818, nc16819, nc16820, nc16821, nc16822, nc16823, nc16824, 
        nc16825, nc16826, nc16827, nc16828, nc16829, 
        \B_DOUT_TEMPR92[39] , \B_DOUT_TEMPR92[38] , 
        \B_DOUT_TEMPR92[37] , \B_DOUT_TEMPR92[36] , 
        \B_DOUT_TEMPR92[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[92][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1644 (.A(\A_DOUT_TEMPR79[6] ), .B(\A_DOUT_TEMPR80[6] ), .C(
        \A_DOUT_TEMPR81[6] ), .D(\A_DOUT_TEMPR82[6] ), .Y(OR4_1644_Y));
    OR4 OR4_2896 (.A(\B_DOUT_TEMPR83[33] ), .B(\B_DOUT_TEMPR84[33] ), 
        .C(\B_DOUT_TEMPR85[33] ), .D(\B_DOUT_TEMPR86[33] ), .Y(
        OR4_2896_Y));
    OR4 OR4_705 (.A(\A_DOUT_TEMPR68[26] ), .B(\A_DOUT_TEMPR69[26] ), 
        .C(\A_DOUT_TEMPR70[26] ), .D(\A_DOUT_TEMPR71[26] ), .Y(
        OR4_705_Y));
    OR2 OR2_74 (.A(\B_DOUT_TEMPR72[15] ), .B(\B_DOUT_TEMPR73[15] ), .Y(
        OR2_74_Y));
    OR4 OR4_1610 (.A(\A_DOUT_TEMPR12[8] ), .B(\A_DOUT_TEMPR13[8] ), .C(
        \A_DOUT_TEMPR14[8] ), .D(\A_DOUT_TEMPR15[8] ), .Y(OR4_1610_Y));
    OR4 OR4_1321 (.A(\B_DOUT_TEMPR87[19] ), .B(\B_DOUT_TEMPR88[19] ), 
        .C(\B_DOUT_TEMPR89[19] ), .D(\B_DOUT_TEMPR90[19] ), .Y(
        OR4_1321_Y));
    OR4 OR4_178 (.A(OR4_327_Y), .B(OR4_2740_Y), .C(OR4_2212_Y), .D(
        OR4_2531_Y), .Y(OR4_178_Y));
    OR4 OR4_634 (.A(OR4_1321_Y), .B(OR4_318_Y), .C(OR4_536_Y), .D(
        OR4_331_Y), .Y(OR4_634_Y));
    OR4 OR4_2463 (.A(\A_DOUT_TEMPR95[36] ), .B(\A_DOUT_TEMPR96[36] ), 
        .C(\A_DOUT_TEMPR97[36] ), .D(\A_DOUT_TEMPR98[36] ), .Y(
        OR4_2463_Y));
    OR4 OR4_1821 (.A(\B_DOUT_TEMPR20[2] ), .B(\B_DOUT_TEMPR21[2] ), .C(
        \B_DOUT_TEMPR22[2] ), .D(\B_DOUT_TEMPR23[2] ), .Y(OR4_1821_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%40%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R40C2 (
        .A_DOUT({nc16830, nc16831, nc16832, nc16833, nc16834, nc16835, 
        nc16836, nc16837, nc16838, nc16839, nc16840, nc16841, nc16842, 
        nc16843, nc16844, \A_DOUT_TEMPR40[14] , \A_DOUT_TEMPR40[13] , 
        \A_DOUT_TEMPR40[12] , \A_DOUT_TEMPR40[11] , 
        \A_DOUT_TEMPR40[10] }), .B_DOUT({nc16845, nc16846, nc16847, 
        nc16848, nc16849, nc16850, nc16851, nc16852, nc16853, nc16854, 
        nc16855, nc16856, nc16857, nc16858, nc16859, 
        \B_DOUT_TEMPR40[14] , \B_DOUT_TEMPR40[13] , 
        \B_DOUT_TEMPR40[12] , \B_DOUT_TEMPR40[11] , 
        \B_DOUT_TEMPR40[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[40][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1018 (.A(\A_DOUT_TEMPR36[25] ), .B(\A_DOUT_TEMPR37[25] ), 
        .C(\A_DOUT_TEMPR38[25] ), .D(\A_DOUT_TEMPR39[25] ), .Y(
        OR4_1018_Y));
    OR4 OR4_2049 (.A(\A_DOUT_TEMPR24[21] ), .B(\A_DOUT_TEMPR25[21] ), 
        .C(\A_DOUT_TEMPR26[21] ), .D(\A_DOUT_TEMPR27[21] ), .Y(
        OR4_2049_Y));
    OR4 OR4_379 (.A(\B_DOUT_TEMPR68[34] ), .B(\B_DOUT_TEMPR69[34] ), 
        .C(\B_DOUT_TEMPR70[34] ), .D(\B_DOUT_TEMPR71[34] ), .Y(
        OR4_379_Y));
    OR4 OR4_392 (.A(OR4_796_Y), .B(OR4_1734_Y), .C(OR4_2201_Y), .D(
        OR4_2991_Y), .Y(OR4_392_Y));
    OR4 OR4_121 (.A(OR4_1_Y), .B(OR4_430_Y), .C(OR4_2673_Y), .D(
        OR4_1587_Y), .Y(OR4_121_Y));
    OR4 OR4_2549 (.A(\A_DOUT_TEMPR8[36] ), .B(\A_DOUT_TEMPR9[36] ), .C(
        \A_DOUT_TEMPR10[36] ), .D(\A_DOUT_TEMPR11[36] ), .Y(OR4_2549_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%54%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R54C4 (
        .A_DOUT({nc16860, nc16861, nc16862, nc16863, nc16864, nc16865, 
        nc16866, nc16867, nc16868, nc16869, nc16870, nc16871, nc16872, 
        nc16873, nc16874, \A_DOUT_TEMPR54[24] , \A_DOUT_TEMPR54[23] , 
        \A_DOUT_TEMPR54[22] , \A_DOUT_TEMPR54[21] , 
        \A_DOUT_TEMPR54[20] }), .B_DOUT({nc16875, nc16876, nc16877, 
        nc16878, nc16879, nc16880, nc16881, nc16882, nc16883, nc16884, 
        nc16885, nc16886, nc16887, nc16888, nc16889, 
        \B_DOUT_TEMPR54[24] , \B_DOUT_TEMPR54[23] , 
        \B_DOUT_TEMPR54[22] , \B_DOUT_TEMPR54[21] , 
        \B_DOUT_TEMPR54[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[54][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%33%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R33C6 (
        .A_DOUT({nc16890, nc16891, nc16892, nc16893, nc16894, nc16895, 
        nc16896, nc16897, nc16898, nc16899, nc16900, nc16901, nc16902, 
        nc16903, nc16904, \A_DOUT_TEMPR33[34] , \A_DOUT_TEMPR33[33] , 
        \A_DOUT_TEMPR33[32] , \A_DOUT_TEMPR33[31] , 
        \A_DOUT_TEMPR33[30] }), .B_DOUT({nc16905, nc16906, nc16907, 
        nc16908, nc16909, nc16910, nc16911, nc16912, nc16913, nc16914, 
        nc16915, nc16916, nc16917, nc16918, nc16919, 
        \B_DOUT_TEMPR33[34] , \B_DOUT_TEMPR33[33] , 
        \B_DOUT_TEMPR33[32] , \B_DOUT_TEMPR33[31] , 
        \B_DOUT_TEMPR33[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[33][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[26]  (.A(OR4_2770_Y), .B(OR4_1629_Y), .C(
        OR4_2309_Y), .D(OR4_660_Y), .Y(B_DOUT[26]));
    OR4 OR4_1276 (.A(OR4_883_Y), .B(OR4_2747_Y), .C(OR4_2278_Y), .D(
        OR4_957_Y), .Y(OR4_1276_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENA[14]  (.A(A_WBYTE_EN[7]), .B(
        A_WEN), .Y(\WBYTEENA[14] ));
    OR4 OR4_2886 (.A(\A_DOUT_TEMPR99[37] ), .B(\A_DOUT_TEMPR100[37] ), 
        .C(\A_DOUT_TEMPR101[37] ), .D(\A_DOUT_TEMPR102[37] ), .Y(
        OR4_2886_Y));
    OR4 OR4_908 (.A(OR4_664_Y), .B(OR4_2746_Y), .C(OR4_2948_Y), .D(
        OR4_2757_Y), .Y(OR4_908_Y));
    OR4 \OR4_A_DOUT[23]  (.A(OR4_2547_Y), .B(OR4_24_Y), .C(OR4_2217_Y), 
        .D(OR4_58_Y), .Y(A_DOUT[23]));
    OR4 OR4_2650 (.A(\B_DOUT_TEMPR87[24] ), .B(\B_DOUT_TEMPR88[24] ), 
        .C(\B_DOUT_TEMPR89[24] ), .D(\B_DOUT_TEMPR90[24] ), .Y(
        OR4_2650_Y));
    OR4 OR4_2342 (.A(\B_DOUT_TEMPR91[33] ), .B(\B_DOUT_TEMPR92[33] ), 
        .C(\B_DOUT_TEMPR93[33] ), .D(\B_DOUT_TEMPR94[33] ), .Y(
        OR4_2342_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%26%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R26C1 (
        .A_DOUT({nc16920, nc16921, nc16922, nc16923, nc16924, nc16925, 
        nc16926, nc16927, nc16928, nc16929, nc16930, nc16931, nc16932, 
        nc16933, nc16934, \A_DOUT_TEMPR26[9] , \A_DOUT_TEMPR26[8] , 
        \A_DOUT_TEMPR26[7] , \A_DOUT_TEMPR26[6] , \A_DOUT_TEMPR26[5] })
        , .B_DOUT({nc16935, nc16936, nc16937, nc16938, nc16939, 
        nc16940, nc16941, nc16942, nc16943, nc16944, nc16945, nc16946, 
        nc16947, nc16948, nc16949, \B_DOUT_TEMPR26[9] , 
        \B_DOUT_TEMPR26[8] , \B_DOUT_TEMPR26[7] , \B_DOUT_TEMPR26[6] , 
        \B_DOUT_TEMPR26[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2790 (.A(\A_DOUT_TEMPR91[26] ), .B(\A_DOUT_TEMPR92[26] ), 
        .C(\A_DOUT_TEMPR93[26] ), .D(\A_DOUT_TEMPR94[26] ), .Y(
        OR4_2790_Y));
    OR4 OR4_2058 (.A(\B_DOUT_TEMPR83[9] ), .B(\B_DOUT_TEMPR84[9] ), .C(
        \B_DOUT_TEMPR85[9] ), .D(\B_DOUT_TEMPR86[9] ), .Y(OR4_2058_Y));
    OR4 OR4_711 (.A(OR4_489_Y), .B(OR4_1313_Y), .C(OR4_361_Y), .D(
        OR4_1287_Y), .Y(OR4_711_Y));
    OR4 OR4_284 (.A(\A_DOUT_TEMPR52[9] ), .B(\A_DOUT_TEMPR53[9] ), .C(
        \A_DOUT_TEMPR54[9] ), .D(\A_DOUT_TEMPR55[9] ), .Y(OR4_284_Y));
    OR4 OR4_272 (.A(\A_DOUT_TEMPR24[15] ), .B(\A_DOUT_TEMPR25[15] ), 
        .C(\A_DOUT_TEMPR26[15] ), .D(\A_DOUT_TEMPR27[15] ), .Y(
        OR4_272_Y));
    OR4 OR4_449 (.A(\B_DOUT_TEMPR64[13] ), .B(\B_DOUT_TEMPR65[13] ), 
        .C(\B_DOUT_TEMPR66[13] ), .D(\B_DOUT_TEMPR67[13] ), .Y(
        OR4_449_Y));
    OR4 OR4_225 (.A(OR4_1822_Y), .B(OR4_2568_Y), .C(OR4_2102_Y), .D(
        OR4_1070_Y), .Y(OR4_225_Y));
    OR4 OR4_595 (.A(\B_DOUT_TEMPR60[11] ), .B(\B_DOUT_TEMPR61[11] ), 
        .C(\B_DOUT_TEMPR62[11] ), .D(\B_DOUT_TEMPR63[11] ), .Y(
        OR4_595_Y));
    OR4 OR4_2516 (.A(\A_DOUT_TEMPR44[24] ), .B(\A_DOUT_TEMPR45[24] ), 
        .C(\A_DOUT_TEMPR46[24] ), .D(\A_DOUT_TEMPR47[24] ), .Y(
        OR4_2516_Y));
    OR4 OR4_108 (.A(\B_DOUT_TEMPR95[27] ), .B(\B_DOUT_TEMPR96[27] ), 
        .C(\B_DOUT_TEMPR97[27] ), .D(\B_DOUT_TEMPR98[27] ), .Y(
        OR4_108_Y));
    OR4 OR4_1114 (.A(\A_DOUT_TEMPR24[32] ), .B(\A_DOUT_TEMPR25[32] ), 
        .C(\A_DOUT_TEMPR26[32] ), .D(\A_DOUT_TEMPR27[32] ), .Y(
        OR4_1114_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%26%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R26C2 (
        .A_DOUT({nc16950, nc16951, nc16952, nc16953, nc16954, nc16955, 
        nc16956, nc16957, nc16958, nc16959, nc16960, nc16961, nc16962, 
        nc16963, nc16964, \A_DOUT_TEMPR26[14] , \A_DOUT_TEMPR26[13] , 
        \A_DOUT_TEMPR26[12] , \A_DOUT_TEMPR26[11] , 
        \A_DOUT_TEMPR26[10] }), .B_DOUT({nc16965, nc16966, nc16967, 
        nc16968, nc16969, nc16970, nc16971, nc16972, nc16973, nc16974, 
        nc16975, nc16976, nc16977, nc16978, nc16979, 
        \B_DOUT_TEMPR26[14] , \B_DOUT_TEMPR26[13] , 
        \B_DOUT_TEMPR26[12] , \B_DOUT_TEMPR26[11] , 
        \B_DOUT_TEMPR26[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_780 (.A(\A_DOUT_TEMPR48[4] ), .B(\A_DOUT_TEMPR49[4] ), .C(
        \A_DOUT_TEMPR50[4] ), .D(\A_DOUT_TEMPR51[4] ), .Y(OR4_780_Y));
    OR4 OR4_2717 (.A(\A_DOUT_TEMPR36[24] ), .B(\A_DOUT_TEMPR37[24] ), 
        .C(\A_DOUT_TEMPR38[24] ), .D(\A_DOUT_TEMPR39[24] ), .Y(
        OR4_2717_Y));
    OR4 OR4_2511 (.A(OR4_1863_Y), .B(OR4_2897_Y), .C(OR4_2325_Y), .D(
        OR4_2726_Y), .Y(OR4_2511_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%20%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R20C6 (
        .A_DOUT({nc16980, nc16981, nc16982, nc16983, nc16984, nc16985, 
        nc16986, nc16987, nc16988, nc16989, nc16990, nc16991, nc16992, 
        nc16993, nc16994, \A_DOUT_TEMPR20[34] , \A_DOUT_TEMPR20[33] , 
        \A_DOUT_TEMPR20[32] , \A_DOUT_TEMPR20[31] , 
        \A_DOUT_TEMPR20[30] }), .B_DOUT({nc16995, nc16996, nc16997, 
        nc16998, nc16999, nc17000, nc17001, nc17002, nc17003, nc17004, 
        nc17005, nc17006, nc17007, nc17008, nc17009, 
        \B_DOUT_TEMPR20[34] , \B_DOUT_TEMPR20[33] , 
        \B_DOUT_TEMPR20[32] , \B_DOUT_TEMPR20[31] , 
        \B_DOUT_TEMPR20[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_309 (.A(\B_DOUT_TEMPR40[24] ), .B(\B_DOUT_TEMPR41[24] ), 
        .C(\B_DOUT_TEMPR42[24] ), .D(\B_DOUT_TEMPR43[24] ), .Y(
        OR4_309_Y));
    OR4 OR4_460 (.A(\A_DOUT_TEMPR111[7] ), .B(\A_DOUT_TEMPR112[7] ), 
        .C(\A_DOUT_TEMPR113[7] ), .D(\A_DOUT_TEMPR114[7] ), .Y(
        OR4_460_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%20%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R20C5 (
        .A_DOUT({nc17010, nc17011, nc17012, nc17013, nc17014, nc17015, 
        nc17016, nc17017, nc17018, nc17019, nc17020, nc17021, nc17022, 
        nc17023, nc17024, \A_DOUT_TEMPR20[29] , \A_DOUT_TEMPR20[28] , 
        \A_DOUT_TEMPR20[27] , \A_DOUT_TEMPR20[26] , 
        \A_DOUT_TEMPR20[25] }), .B_DOUT({nc17025, nc17026, nc17027, 
        nc17028, nc17029, nc17030, nc17031, nc17032, nc17033, nc17034, 
        nc17035, nc17036, nc17037, nc17038, nc17039, 
        \B_DOUT_TEMPR20[29] , \B_DOUT_TEMPR20[28] , 
        \B_DOUT_TEMPR20[27] , \B_DOUT_TEMPR20[26] , 
        \B_DOUT_TEMPR20[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_61 (.A(\B_DOUT_TEMPR72[24] ), .B(\B_DOUT_TEMPR73[24] ), .Y(
        OR2_61_Y));
    OR4 OR4_626 (.A(\B_DOUT_TEMPR115[13] ), .B(\B_DOUT_TEMPR116[13] ), 
        .C(\B_DOUT_TEMPR117[13] ), .D(\B_DOUT_TEMPR118[13] ), .Y(
        OR4_626_Y));
    OR4 OR4_1809 (.A(\B_DOUT_TEMPR56[31] ), .B(\B_DOUT_TEMPR57[31] ), 
        .C(\B_DOUT_TEMPR58[31] ), .D(\B_DOUT_TEMPR59[31] ), .Y(
        OR4_1809_Y));
    OR4 OR4_2780 (.A(\B_DOUT_TEMPR36[13] ), .B(\B_DOUT_TEMPR37[13] ), 
        .C(\B_DOUT_TEMPR38[13] ), .D(\B_DOUT_TEMPR39[13] ), .Y(
        OR4_2780_Y));
    OR4 OR4_2545 (.A(\B_DOUT_TEMPR52[2] ), .B(\B_DOUT_TEMPR53[2] ), .C(
        \B_DOUT_TEMPR54[2] ), .D(\B_DOUT_TEMPR55[2] ), .Y(OR4_2545_Y));
    OR4 OR4_1876 (.A(\A_DOUT_TEMPR64[35] ), .B(\A_DOUT_TEMPR65[35] ), 
        .C(\A_DOUT_TEMPR66[35] ), .D(\A_DOUT_TEMPR67[35] ), .Y(
        OR4_1876_Y));
    OR4 OR4_812 (.A(\B_DOUT_TEMPR52[36] ), .B(\B_DOUT_TEMPR53[36] ), 
        .C(\B_DOUT_TEMPR54[36] ), .D(\B_DOUT_TEMPR55[36] ), .Y(
        OR4_812_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%105%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R105C5 (
        .A_DOUT({nc17040, nc17041, nc17042, nc17043, nc17044, nc17045, 
        nc17046, nc17047, nc17048, nc17049, nc17050, nc17051, nc17052, 
        nc17053, nc17054, \A_DOUT_TEMPR105[29] , \A_DOUT_TEMPR105[28] , 
        \A_DOUT_TEMPR105[27] , \A_DOUT_TEMPR105[26] , 
        \A_DOUT_TEMPR105[25] }), .B_DOUT({nc17055, nc17056, nc17057, 
        nc17058, nc17059, nc17060, nc17061, nc17062, nc17063, nc17064, 
        nc17065, nc17066, nc17067, nc17068, nc17069, 
        \B_DOUT_TEMPR105[29] , \B_DOUT_TEMPR105[28] , 
        \B_DOUT_TEMPR105[27] , \B_DOUT_TEMPR105[26] , 
        \B_DOUT_TEMPR105[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[105][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%73%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R73C4 (
        .A_DOUT({nc17070, nc17071, nc17072, nc17073, nc17074, nc17075, 
        nc17076, nc17077, nc17078, nc17079, nc17080, nc17081, nc17082, 
        nc17083, nc17084, \A_DOUT_TEMPR73[24] , \A_DOUT_TEMPR73[23] , 
        \A_DOUT_TEMPR73[22] , \A_DOUT_TEMPR73[21] , 
        \A_DOUT_TEMPR73[20] }), .B_DOUT({nc17085, nc17086, nc17087, 
        nc17088, nc17089, nc17090, nc17091, nc17092, nc17093, nc17094, 
        nc17095, nc17096, nc17097, nc17098, nc17099, 
        \B_DOUT_TEMPR73[24] , \B_DOUT_TEMPR73[23] , 
        \B_DOUT_TEMPR73[22] , \B_DOUT_TEMPR73[21] , 
        \B_DOUT_TEMPR73[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[73][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_11 (.A(\A_DOUT_TEMPR72[14] ), .B(\A_DOUT_TEMPR73[14] ), .Y(
        OR2_11_Y));
    OR4 OR4_2178 (.A(\A_DOUT_TEMPR75[39] ), .B(\A_DOUT_TEMPR76[39] ), 
        .C(\A_DOUT_TEMPR77[39] ), .D(\A_DOUT_TEMPR78[39] ), .Y(
        OR4_2178_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%34%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R34C4 (
        .A_DOUT({nc17100, nc17101, nc17102, nc17103, nc17104, nc17105, 
        nc17106, nc17107, nc17108, nc17109, nc17110, nc17111, nc17112, 
        nc17113, nc17114, \A_DOUT_TEMPR34[24] , \A_DOUT_TEMPR34[23] , 
        \A_DOUT_TEMPR34[22] , \A_DOUT_TEMPR34[21] , 
        \A_DOUT_TEMPR34[20] }), .B_DOUT({nc17115, nc17116, nc17117, 
        nc17118, nc17119, nc17120, nc17121, nc17122, nc17123, nc17124, 
        nc17125, nc17126, nc17127, nc17128, nc17129, 
        \B_DOUT_TEMPR34[24] , \B_DOUT_TEMPR34[23] , 
        \B_DOUT_TEMPR34[22] , \B_DOUT_TEMPR34[21] , 
        \B_DOUT_TEMPR34[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[34][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_0 (.A(\A_DOUT_TEMPR72[27] ), .B(\A_DOUT_TEMPR73[27] ), .Y(
        OR2_0_Y));
    OR4 OR4_141 (.A(\B_DOUT_TEMPR75[23] ), .B(\B_DOUT_TEMPR76[23] ), 
        .C(\B_DOUT_TEMPR77[23] ), .D(\B_DOUT_TEMPR78[23] ), .Y(
        OR4_141_Y));
    OR4 OR4_2397 (.A(\B_DOUT_TEMPR44[16] ), .B(\B_DOUT_TEMPR45[16] ), 
        .C(\B_DOUT_TEMPR46[16] ), .D(\B_DOUT_TEMPR47[16] ), .Y(
        OR4_2397_Y));
    OR4 OR4_2292 (.A(\A_DOUT_TEMPR8[6] ), .B(\A_DOUT_TEMPR9[6] ), .C(
        \A_DOUT_TEMPR10[6] ), .D(\A_DOUT_TEMPR11[6] ), .Y(OR4_2292_Y));
    OR4 OR4_358 (.A(\B_DOUT_TEMPR36[38] ), .B(\B_DOUT_TEMPR37[38] ), 
        .C(\B_DOUT_TEMPR38[38] ), .D(\B_DOUT_TEMPR39[38] ), .Y(
        OR4_358_Y));
    OR4 OR4_1101 (.A(OR4_1656_Y), .B(OR4_1017_Y), .C(OR2_75_Y), .D(
        \B_DOUT_TEMPR74[8] ), .Y(OR4_1101_Y));
    OR4 OR4_637 (.A(\B_DOUT_TEMPR56[1] ), .B(\B_DOUT_TEMPR57[1] ), .C(
        \B_DOUT_TEMPR58[1] ), .D(\B_DOUT_TEMPR59[1] ), .Y(OR4_637_Y));
    OR4 OR4_2154 (.A(\B_DOUT_TEMPR0[18] ), .B(\B_DOUT_TEMPR1[18] ), .C(
        \B_DOUT_TEMPR2[18] ), .D(\B_DOUT_TEMPR3[18] ), .Y(OR4_2154_Y));
    OR4 OR4_755 (.A(\A_DOUT_TEMPR60[1] ), .B(\A_DOUT_TEMPR61[1] ), .C(
        \A_DOUT_TEMPR62[1] ), .D(\A_DOUT_TEMPR63[1] ), .Y(OR4_755_Y));
    OR4 OR4_1815 (.A(\B_DOUT_TEMPR52[24] ), .B(\B_DOUT_TEMPR53[24] ), 
        .C(\B_DOUT_TEMPR54[24] ), .D(\B_DOUT_TEMPR55[24] ), .Y(
        OR4_1815_Y));
    OR4 OR4_1640 (.A(OR4_2598_Y), .B(OR4_356_Y), .C(OR2_61_Y), .D(
        \B_DOUT_TEMPR74[24] ), .Y(OR4_1640_Y));
    OR4 OR4_202 (.A(\B_DOUT_TEMPR87[4] ), .B(\B_DOUT_TEMPR88[4] ), .C(
        \B_DOUT_TEMPR89[4] ), .D(\B_DOUT_TEMPR90[4] ), .Y(OR4_202_Y));
    OR4 OR4_2873 (.A(OR4_3008_Y), .B(OR4_254_Y), .C(OR4_2951_Y), .D(
        OR4_269_Y), .Y(OR4_2873_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%11%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R11C0 (
        .A_DOUT({nc17130, nc17131, nc17132, nc17133, nc17134, nc17135, 
        nc17136, nc17137, nc17138, nc17139, nc17140, nc17141, nc17142, 
        nc17143, nc17144, \A_DOUT_TEMPR11[4] , \A_DOUT_TEMPR11[3] , 
        \A_DOUT_TEMPR11[2] , \A_DOUT_TEMPR11[1] , \A_DOUT_TEMPR11[0] })
        , .B_DOUT({nc17145, nc17146, nc17147, nc17148, nc17149, 
        nc17150, nc17151, nc17152, nc17153, nc17154, nc17155, nc17156, 
        nc17157, nc17158, nc17159, \B_DOUT_TEMPR11[4] , 
        \B_DOUT_TEMPR11[3] , \B_DOUT_TEMPR11[2] , \B_DOUT_TEMPR11[1] , 
        \B_DOUT_TEMPR11[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1005 (.A(\A_DOUT_TEMPR4[37] ), .B(\A_DOUT_TEMPR5[37] ), .C(
        \A_DOUT_TEMPR6[37] ), .D(\A_DOUT_TEMPR7[37] ), .Y(OR4_1005_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[12]  (.A(CFG3_12_Y), .B(
        CFG3_15_Y), .Y(\BLKY2[12] ));
    OR4 OR4_2931 (.A(\A_DOUT_TEMPR99[31] ), .B(\A_DOUT_TEMPR100[31] ), 
        .C(\A_DOUT_TEMPR101[31] ), .D(\A_DOUT_TEMPR102[31] ), .Y(
        OR4_2931_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%44%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R44C6 (
        .A_DOUT({nc17160, nc17161, nc17162, nc17163, nc17164, nc17165, 
        nc17166, nc17167, nc17168, nc17169, nc17170, nc17171, nc17172, 
        nc17173, nc17174, \A_DOUT_TEMPR44[34] , \A_DOUT_TEMPR44[33] , 
        \A_DOUT_TEMPR44[32] , \A_DOUT_TEMPR44[31] , 
        \A_DOUT_TEMPR44[30] }), .B_DOUT({nc17175, nc17176, nc17177, 
        nc17178, nc17179, nc17180, nc17181, nc17182, nc17183, nc17184, 
        nc17185, nc17186, nc17187, nc17188, nc17189, 
        \B_DOUT_TEMPR44[34] , \B_DOUT_TEMPR44[33] , 
        \B_DOUT_TEMPR44[32] , \B_DOUT_TEMPR44[31] , 
        \B_DOUT_TEMPR44[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[44][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1158 (.A(OR4_197_Y), .B(OR4_1491_Y), .C(OR4_1237_Y), .D(
        OR4_1828_Y), .Y(OR4_1158_Y));
    OR4 OR4_1048 (.A(\A_DOUT_TEMPR60[0] ), .B(\A_DOUT_TEMPR61[0] ), .C(
        \A_DOUT_TEMPR62[0] ), .D(\A_DOUT_TEMPR63[0] ), .Y(OR4_1048_Y));
    OR4 OR4_2266 (.A(OR4_1804_Y), .B(OR4_2633_Y), .C(OR4_1676_Y), .D(
        OR4_1818_Y), .Y(OR4_2266_Y));
    OR4 OR4_124 (.A(\B_DOUT_TEMPR64[18] ), .B(\B_DOUT_TEMPR65[18] ), 
        .C(\B_DOUT_TEMPR66[18] ), .D(\B_DOUT_TEMPR67[18] ), .Y(
        OR4_124_Y));
    OR4 OR4_1931 (.A(\A_DOUT_TEMPR20[17] ), .B(\A_DOUT_TEMPR21[17] ), 
        .C(\A_DOUT_TEMPR22[17] ), .D(\A_DOUT_TEMPR23[17] ), .Y(
        OR4_1931_Y));
    OR4 OR4_324 (.A(OR4_2644_Y), .B(OR4_2952_Y), .C(OR4_1489_Y), .D(
        OR4_2399_Y), .Y(OR4_324_Y));
    OR4 OR4_2779 (.A(\B_DOUT_TEMPR115[6] ), .B(\B_DOUT_TEMPR116[6] ), 
        .C(\B_DOUT_TEMPR117[6] ), .D(\B_DOUT_TEMPR118[6] ), .Y(
        OR4_2779_Y));
    OR4 OR4_2494 (.A(\B_DOUT_TEMPR111[18] ), .B(\B_DOUT_TEMPR112[18] ), 
        .C(\B_DOUT_TEMPR113[18] ), .D(\B_DOUT_TEMPR114[18] ), .Y(
        OR4_2494_Y));
    OR4 OR4_2387 (.A(\B_DOUT_TEMPR87[14] ), .B(\B_DOUT_TEMPR88[14] ), 
        .C(\B_DOUT_TEMPR89[14] ), .D(\B_DOUT_TEMPR90[14] ), .Y(
        OR4_2387_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%67%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R67C4 (
        .A_DOUT({nc17190, nc17191, nc17192, nc17193, nc17194, nc17195, 
        nc17196, nc17197, nc17198, nc17199, nc17200, nc17201, nc17202, 
        nc17203, nc17204, \A_DOUT_TEMPR67[24] , \A_DOUT_TEMPR67[23] , 
        \A_DOUT_TEMPR67[22] , \A_DOUT_TEMPR67[21] , 
        \A_DOUT_TEMPR67[20] }), .B_DOUT({nc17205, nc17206, nc17207, 
        nc17208, nc17209, nc17210, nc17211, nc17212, nc17213, nc17214, 
        nc17215, nc17216, nc17217, nc17218, nc17219, 
        \B_DOUT_TEMPR67[24] , \B_DOUT_TEMPR67[23] , 
        \B_DOUT_TEMPR67[22] , \B_DOUT_TEMPR67[21] , 
        \B_DOUT_TEMPR67[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[67][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_169 (.A(\B_DOUT_TEMPR8[25] ), .B(\B_DOUT_TEMPR9[25] ), .C(
        \B_DOUT_TEMPR10[25] ), .D(\B_DOUT_TEMPR11[25] ), .Y(OR4_169_Y));
    OR4 OR4_2282 (.A(\B_DOUT_TEMPR16[20] ), .B(\B_DOUT_TEMPR17[20] ), 
        .C(\B_DOUT_TEMPR18[20] ), .D(\B_DOUT_TEMPR19[20] ), .Y(
        OR4_2282_Y));
    OR4 OR4_2948 (.A(\B_DOUT_TEMPR95[11] ), .B(\B_DOUT_TEMPR96[11] ), 
        .C(\B_DOUT_TEMPR97[11] ), .D(\B_DOUT_TEMPR98[11] ), .Y(
        OR4_2948_Y));
    OR4 OR4_1770 (.A(\B_DOUT_TEMPR111[2] ), .B(\B_DOUT_TEMPR112[2] ), 
        .C(\B_DOUT_TEMPR113[2] ), .D(\B_DOUT_TEMPR114[2] ), .Y(
        OR4_1770_Y));
    OR4 OR4_245 (.A(\A_DOUT_TEMPR79[8] ), .B(\A_DOUT_TEMPR80[8] ), .C(
        \A_DOUT_TEMPR81[8] ), .D(\A_DOUT_TEMPR82[8] ), .Y(OR4_245_Y));
    OR4 OR4_958 (.A(\A_DOUT_TEMPR99[36] ), .B(\A_DOUT_TEMPR100[36] ), 
        .C(\A_DOUT_TEMPR101[36] ), .D(\A_DOUT_TEMPR102[36] ), .Y(
        OR4_958_Y));
    OR4 OR4_1853 (.A(OR4_2997_Y), .B(OR4_1089_Y), .C(OR4_237_Y), .D(
        OR4_2194_Y), .Y(OR4_1853_Y));
    OR4 OR4_1927 (.A(\B_DOUT_TEMPR95[23] ), .B(\B_DOUT_TEMPR96[23] ), 
        .C(\B_DOUT_TEMPR97[23] ), .D(\B_DOUT_TEMPR98[23] ), .Y(
        OR4_1927_Y));
    OR4 OR4_2855 (.A(\B_DOUT_TEMPR44[21] ), .B(\B_DOUT_TEMPR45[21] ), 
        .C(\B_DOUT_TEMPR46[21] ), .D(\B_DOUT_TEMPR47[21] ), .Y(
        OR4_2855_Y));
    OR4 OR4_1807 (.A(\B_DOUT_TEMPR111[26] ), .B(\B_DOUT_TEMPR112[26] ), 
        .C(\B_DOUT_TEMPR113[26] ), .D(\B_DOUT_TEMPR114[26] ), .Y(
        OR4_1807_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%2%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R2C6 (
        .A_DOUT({nc17220, nc17221, nc17222, nc17223, nc17224, nc17225, 
        nc17226, nc17227, nc17228, nc17229, nc17230, nc17231, nc17232, 
        nc17233, nc17234, \A_DOUT_TEMPR2[34] , \A_DOUT_TEMPR2[33] , 
        \A_DOUT_TEMPR2[32] , \A_DOUT_TEMPR2[31] , \A_DOUT_TEMPR2[30] })
        , .B_DOUT({nc17235, nc17236, nc17237, nc17238, nc17239, 
        nc17240, nc17241, nc17242, nc17243, nc17244, nc17245, nc17246, 
        nc17247, nc17248, nc17249, \B_DOUT_TEMPR2[34] , 
        \B_DOUT_TEMPR2[33] , \B_DOUT_TEMPR2[32] , \B_DOUT_TEMPR2[31] , 
        \B_DOUT_TEMPR2[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%71%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R71C4 (
        .A_DOUT({nc17250, nc17251, nc17252, nc17253, nc17254, nc17255, 
        nc17256, nc17257, nc17258, nc17259, nc17260, nc17261, nc17262, 
        nc17263, nc17264, \A_DOUT_TEMPR71[24] , \A_DOUT_TEMPR71[23] , 
        \A_DOUT_TEMPR71[22] , \A_DOUT_TEMPR71[21] , 
        \A_DOUT_TEMPR71[20] }), .B_DOUT({nc17265, nc17266, nc17267, 
        nc17268, nc17269, nc17270, nc17271, nc17272, nc17273, nc17274, 
        nc17275, nc17276, nc17277, nc17278, nc17279, 
        \B_DOUT_TEMPR71[24] , \B_DOUT_TEMPR71[23] , 
        \B_DOUT_TEMPR71[22] , \B_DOUT_TEMPR71[21] , 
        \B_DOUT_TEMPR71[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[71][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2176 (.A(\B_DOUT_TEMPR4[5] ), .B(\B_DOUT_TEMPR5[5] ), .C(
        \B_DOUT_TEMPR6[5] ), .D(\B_DOUT_TEMPR7[5] ), .Y(OR4_2176_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%108%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R108C7 (
        .A_DOUT({nc17280, nc17281, nc17282, nc17283, nc17284, nc17285, 
        nc17286, nc17287, nc17288, nc17289, nc17290, nc17291, nc17292, 
        nc17293, nc17294, \A_DOUT_TEMPR108[39] , \A_DOUT_TEMPR108[38] , 
        \A_DOUT_TEMPR108[37] , \A_DOUT_TEMPR108[36] , 
        \A_DOUT_TEMPR108[35] }), .B_DOUT({nc17295, nc17296, nc17297, 
        nc17298, nc17299, nc17300, nc17301, nc17302, nc17303, nc17304, 
        nc17305, nc17306, nc17307, nc17308, nc17309, 
        \B_DOUT_TEMPR108[39] , \B_DOUT_TEMPR108[38] , 
        \B_DOUT_TEMPR108[37] , \B_DOUT_TEMPR108[36] , 
        \B_DOUT_TEMPR108[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[108][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2578 (.A(\B_DOUT_TEMPR44[29] ), .B(\B_DOUT_TEMPR45[29] ), 
        .C(\B_DOUT_TEMPR46[29] ), .D(\B_DOUT_TEMPR47[29] ), .Y(
        OR4_2578_Y));
    OR4 OR4_237 (.A(\B_DOUT_TEMPR79[1] ), .B(\B_DOUT_TEMPR80[1] ), .C(
        \B_DOUT_TEMPR81[1] ), .D(\B_DOUT_TEMPR82[1] ), .Y(OR4_237_Y));
    OR4 OR4_646 (.A(OR4_218_Y), .B(OR4_2176_Y), .C(OR4_822_Y), .D(
        OR4_1799_Y), .Y(OR4_646_Y));
    OR4 OR4_1759 (.A(OR4_2145_Y), .B(OR4_805_Y), .C(OR4_2153_Y), .D(
        OR4_2445_Y), .Y(OR4_1759_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%63%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R63C6 (
        .A_DOUT({nc17310, nc17311, nc17312, nc17313, nc17314, nc17315, 
        nc17316, nc17317, nc17318, nc17319, nc17320, nc17321, nc17322, 
        nc17323, nc17324, \A_DOUT_TEMPR63[34] , \A_DOUT_TEMPR63[33] , 
        \A_DOUT_TEMPR63[32] , \A_DOUT_TEMPR63[31] , 
        \A_DOUT_TEMPR63[30] }), .B_DOUT({nc17325, nc17326, nc17327, 
        nc17328, nc17329, nc17330, nc17331, nc17332, nc17333, nc17334, 
        nc17335, nc17336, nc17337, nc17338, nc17339, 
        \B_DOUT_TEMPR63[34] , \B_DOUT_TEMPR63[33] , 
        \B_DOUT_TEMPR63[32] , \B_DOUT_TEMPR63[31] , 
        \B_DOUT_TEMPR63[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[63][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%52%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R52C7 (
        .A_DOUT({nc17340, nc17341, nc17342, nc17343, nc17344, nc17345, 
        nc17346, nc17347, nc17348, nc17349, nc17350, nc17351, nc17352, 
        nc17353, nc17354, \A_DOUT_TEMPR52[39] , \A_DOUT_TEMPR52[38] , 
        \A_DOUT_TEMPR52[37] , \A_DOUT_TEMPR52[36] , 
        \A_DOUT_TEMPR52[35] }), .B_DOUT({nc17355, nc17356, nc17357, 
        nc17358, nc17359, nc17360, nc17361, nc17362, nc17363, nc17364, 
        nc17365, nc17366, nc17367, nc17368, nc17369, 
        \B_DOUT_TEMPR52[39] , \B_DOUT_TEMPR52[38] , 
        \B_DOUT_TEMPR52[37] , \B_DOUT_TEMPR52[36] , 
        \B_DOUT_TEMPR52[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[52][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%28%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R28C5 (
        .A_DOUT({nc17370, nc17371, nc17372, nc17373, nc17374, nc17375, 
        nc17376, nc17377, nc17378, nc17379, nc17380, nc17381, nc17382, 
        nc17383, nc17384, \A_DOUT_TEMPR28[29] , \A_DOUT_TEMPR28[28] , 
        \A_DOUT_TEMPR28[27] , \A_DOUT_TEMPR28[26] , 
        \A_DOUT_TEMPR28[25] }), .B_DOUT({nc17385, nc17386, nc17387, 
        nc17388, nc17389, nc17390, nc17391, nc17392, nc17393, nc17394, 
        nc17395, nc17396, nc17397, nc17398, nc17399, 
        \B_DOUT_TEMPR28[29] , \B_DOUT_TEMPR28[28] , 
        \B_DOUT_TEMPR28[27] , \B_DOUT_TEMPR28[26] , 
        \B_DOUT_TEMPR28[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[18]  (.A(OR4_2752_Y), .B(OR4_877_Y), .C(OR4_2609_Y)
        , .D(OR4_1430_Y), .Y(B_DOUT[18]));
    OR4 OR4_2605 (.A(\B_DOUT_TEMPR103[10] ), .B(\B_DOUT_TEMPR104[10] ), 
        .C(\B_DOUT_TEMPR105[10] ), .D(\B_DOUT_TEMPR106[10] ), .Y(
        OR4_2605_Y));
    OR4 OR4_2233 (.A(\A_DOUT_TEMPR8[4] ), .B(\A_DOUT_TEMPR9[4] ), .C(
        \A_DOUT_TEMPR10[4] ), .D(\A_DOUT_TEMPR11[4] ), .Y(OR4_2233_Y));
    OR4 OR4_2484 (.A(OR4_2499_Y), .B(OR4_2761_Y), .C(OR4_1203_Y), .D(
        OR4_2763_Y), .Y(OR4_2484_Y));
    OR4 OR4_158 (.A(\B_DOUT_TEMPR20[33] ), .B(\B_DOUT_TEMPR21[33] ), 
        .C(\B_DOUT_TEMPR22[33] ), .D(\B_DOUT_TEMPR23[33] ), .Y(
        OR4_158_Y));
    OR4 OR4_1233 (.A(\B_DOUT_TEMPR103[19] ), .B(\B_DOUT_TEMPR104[19] ), 
        .C(\B_DOUT_TEMPR105[19] ), .D(\B_DOUT_TEMPR106[19] ), .Y(
        OR4_1233_Y));
    OR4 OR4_1144 (.A(\B_DOUT_TEMPR32[25] ), .B(\B_DOUT_TEMPR33[25] ), 
        .C(\B_DOUT_TEMPR34[25] ), .D(\B_DOUT_TEMPR35[25] ), .Y(
        OR4_1144_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%115%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R115C0 (
        .A_DOUT({nc17400, nc17401, nc17402, nc17403, nc17404, nc17405, 
        nc17406, nc17407, nc17408, nc17409, nc17410, nc17411, nc17412, 
        nc17413, nc17414, \A_DOUT_TEMPR115[4] , \A_DOUT_TEMPR115[3] , 
        \A_DOUT_TEMPR115[2] , \A_DOUT_TEMPR115[1] , 
        \A_DOUT_TEMPR115[0] }), .B_DOUT({nc17415, nc17416, nc17417, 
        nc17418, nc17419, nc17420, nc17421, nc17422, nc17423, nc17424, 
        nc17425, nc17426, nc17427, nc17428, nc17429, 
        \B_DOUT_TEMPR115[4] , \B_DOUT_TEMPR115[3] , 
        \B_DOUT_TEMPR115[2] , \B_DOUT_TEMPR115[1] , 
        \B_DOUT_TEMPR115[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[115][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%116%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R116C4 (
        .A_DOUT({nc17430, nc17431, nc17432, nc17433, nc17434, nc17435, 
        nc17436, nc17437, nc17438, nc17439, nc17440, nc17441, nc17442, 
        nc17443, nc17444, \A_DOUT_TEMPR116[24] , \A_DOUT_TEMPR116[23] , 
        \A_DOUT_TEMPR116[22] , \A_DOUT_TEMPR116[21] , 
        \A_DOUT_TEMPR116[20] }), .B_DOUT({nc17445, nc17446, nc17447, 
        nc17448, nc17449, nc17450, nc17451, nc17452, nc17453, nc17454, 
        nc17455, nc17456, nc17457, nc17458, nc17459, 
        \B_DOUT_TEMPR116[24] , \B_DOUT_TEMPR116[23] , 
        \B_DOUT_TEMPR116[22] , \B_DOUT_TEMPR116[21] , 
        \B_DOUT_TEMPR116[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[116][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_359 (.A(\A_DOUT_TEMPR24[34] ), .B(\A_DOUT_TEMPR25[34] ), 
        .C(\A_DOUT_TEMPR26[34] ), .D(\A_DOUT_TEMPR27[34] ), .Y(
        OR4_359_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%71%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R71C3 (
        .A_DOUT({nc17460, nc17461, nc17462, nc17463, nc17464, nc17465, 
        nc17466, nc17467, nc17468, nc17469, nc17470, nc17471, nc17472, 
        nc17473, nc17474, \A_DOUT_TEMPR71[19] , \A_DOUT_TEMPR71[18] , 
        \A_DOUT_TEMPR71[17] , \A_DOUT_TEMPR71[16] , 
        \A_DOUT_TEMPR71[15] }), .B_DOUT({nc17475, nc17476, nc17477, 
        nc17478, nc17479, nc17480, nc17481, nc17482, nc17483, nc17484, 
        nc17485, nc17486, nc17487, nc17488, nc17489, 
        \B_DOUT_TEMPR71[19] , \B_DOUT_TEMPR71[18] , 
        \B_DOUT_TEMPR71[17] , \B_DOUT_TEMPR71[16] , 
        \B_DOUT_TEMPR71[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[71][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1156 (.A(\A_DOUT_TEMPR0[4] ), .B(\A_DOUT_TEMPR1[4] ), .C(
        \A_DOUT_TEMPR2[4] ), .D(\A_DOUT_TEMPR3[4] ), .Y(OR4_1156_Y));
    OR4 OR4_932 (.A(\B_DOUT_TEMPR83[13] ), .B(\B_DOUT_TEMPR84[13] ), 
        .C(\B_DOUT_TEMPR85[13] ), .D(\B_DOUT_TEMPR86[13] ), .Y(
        OR4_932_Y));
    OR4 OR4_2866 (.A(\A_DOUT_TEMPR28[19] ), .B(\A_DOUT_TEMPR29[19] ), 
        .C(\A_DOUT_TEMPR30[19] ), .D(\A_DOUT_TEMPR31[19] ), .Y(
        OR4_2866_Y));
    OR4 OR4_1593 (.A(\B_DOUT_TEMPR111[9] ), .B(\B_DOUT_TEMPR112[9] ), 
        .C(\B_DOUT_TEMPR113[9] ), .D(\B_DOUT_TEMPR114[9] ), .Y(
        OR4_1593_Y));
    OR4 OR4_1377 (.A(\A_DOUT_TEMPR40[30] ), .B(\A_DOUT_TEMPR41[30] ), 
        .C(\A_DOUT_TEMPR42[30] ), .D(\A_DOUT_TEMPR43[30] ), .Y(
        OR4_1377_Y));
    OR4 OR4_1558 (.A(\A_DOUT_TEMPR111[14] ), .B(\A_DOUT_TEMPR112[14] ), 
        .C(\A_DOUT_TEMPR113[14] ), .D(\A_DOUT_TEMPR114[14] ), .Y(
        OR4_1558_Y));
    OR4 OR4_1820 (.A(\B_DOUT_TEMPR24[7] ), .B(\B_DOUT_TEMPR25[7] ), .C(
        \B_DOUT_TEMPR26[7] ), .D(\B_DOUT_TEMPR27[7] ), .Y(OR4_1820_Y));
    OR4 OR4_135 (.A(OR4_112_Y), .B(OR4_508_Y), .C(OR4_1267_Y), .D(
        OR4_2067_Y), .Y(OR4_135_Y));
    OR4 OR4_1272 (.A(\A_DOUT_TEMPR16[8] ), .B(\A_DOUT_TEMPR17[8] ), .C(
        \A_DOUT_TEMPR18[8] ), .D(\A_DOUT_TEMPR19[8] ), .Y(OR4_1272_Y));
    OR4 OR4_2147 (.A(\A_DOUT_TEMPR28[14] ), .B(\A_DOUT_TEMPR29[14] ), 
        .C(\A_DOUT_TEMPR30[14] ), .D(\A_DOUT_TEMPR31[14] ), .Y(
        OR4_2147_Y));
    OR4 OR4_717 (.A(\B_DOUT_TEMPR36[11] ), .B(\B_DOUT_TEMPR37[11] ), 
        .C(\B_DOUT_TEMPR38[11] ), .D(\B_DOUT_TEMPR39[11] ), .Y(
        OR4_717_Y));
    OR4 OR4_2644 (.A(\A_DOUT_TEMPR0[32] ), .B(\A_DOUT_TEMPR1[32] ), .C(
        \A_DOUT_TEMPR2[32] ), .D(\A_DOUT_TEMPR3[32] ), .Y(OR4_2644_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%21%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R21C7 (
        .A_DOUT({nc17490, nc17491, nc17492, nc17493, nc17494, nc17495, 
        nc17496, nc17497, nc17498, nc17499, nc17500, nc17501, nc17502, 
        nc17503, nc17504, \A_DOUT_TEMPR21[39] , \A_DOUT_TEMPR21[38] , 
        \A_DOUT_TEMPR21[37] , \A_DOUT_TEMPR21[36] , 
        \A_DOUT_TEMPR21[35] }), .B_DOUT({nc17505, nc17506, nc17507, 
        nc17508, nc17509, nc17510, nc17511, nc17512, nc17513, nc17514, 
        nc17515, nc17516, nc17517, nc17518, nc17519, 
        \B_DOUT_TEMPR21[39] , \B_DOUT_TEMPR21[38] , 
        \B_DOUT_TEMPR21[37] , \B_DOUT_TEMPR21[36] , 
        \B_DOUT_TEMPR21[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1193 (.A(\A_DOUT_TEMPR99[34] ), .B(\A_DOUT_TEMPR100[34] ), 
        .C(\A_DOUT_TEMPR101[34] ), .D(\A_DOUT_TEMPR102[34] ), .Y(
        OR4_1193_Y));
    OR4 OR4_313 (.A(OR4_188_Y), .B(OR4_1871_Y), .C(OR4_1327_Y), .D(
        OR4_2639_Y), .Y(OR4_313_Y));
    OR4 OR4_930 (.A(\B_DOUT_TEMPR8[17] ), .B(\B_DOUT_TEMPR9[17] ), .C(
        \B_DOUT_TEMPR10[17] ), .D(\B_DOUT_TEMPR11[17] ), .Y(OR4_930_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%113%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R113C3 (
        .A_DOUT({nc17520, nc17521, nc17522, nc17523, nc17524, nc17525, 
        nc17526, nc17527, nc17528, nc17529, nc17530, nc17531, nc17532, 
        nc17533, nc17534, \A_DOUT_TEMPR113[19] , \A_DOUT_TEMPR113[18] , 
        \A_DOUT_TEMPR113[17] , \A_DOUT_TEMPR113[16] , 
        \A_DOUT_TEMPR113[15] }), .B_DOUT({nc17535, nc17536, nc17537, 
        nc17538, nc17539, nc17540, nc17541, nc17542, nc17543, nc17544, 
        nc17545, nc17546, nc17547, nc17548, nc17549, 
        \B_DOUT_TEMPR113[19] , \B_DOUT_TEMPR113[18] , 
        \B_DOUT_TEMPR113[17] , \B_DOUT_TEMPR113[16] , 
        \B_DOUT_TEMPR113[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[113][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_761 (.A(\A_DOUT_TEMPR40[13] ), .B(\A_DOUT_TEMPR41[13] ), 
        .C(\A_DOUT_TEMPR42[13] ), .D(\A_DOUT_TEMPR43[13] ), .Y(
        OR4_761_Y));
    OR4 OR4_2607 (.A(\A_DOUT_TEMPR32[0] ), .B(\A_DOUT_TEMPR33[0] ), .C(
        \A_DOUT_TEMPR34[0] ), .D(\A_DOUT_TEMPR35[0] ), .Y(OR4_2607_Y));
    OR4 OR4_718 (.A(\A_DOUT_TEMPR103[24] ), .B(\A_DOUT_TEMPR104[24] ), 
        .C(\A_DOUT_TEMPR105[24] ), .D(\A_DOUT_TEMPR106[24] ), .Y(
        OR4_718_Y));
    OR4 OR4_1824 (.A(\B_DOUT_TEMPR68[15] ), .B(\B_DOUT_TEMPR69[15] ), 
        .C(\B_DOUT_TEMPR70[15] ), .D(\B_DOUT_TEMPR71[15] ), .Y(
        OR4_1824_Y));
    OR4 OR4_1092 (.A(\A_DOUT_TEMPR8[14] ), .B(\A_DOUT_TEMPR9[14] ), .C(
        \A_DOUT_TEMPR10[14] ), .D(\A_DOUT_TEMPR11[14] ), .Y(OR4_1092_Y)
        );
    OR4 OR4_2294 (.A(\B_DOUT_TEMPR99[23] ), .B(\B_DOUT_TEMPR100[23] ), 
        .C(\B_DOUT_TEMPR101[23] ), .D(\B_DOUT_TEMPR102[23] ), .Y(
        OR4_2294_Y));
    OR4 OR4_613 (.A(\A_DOUT_TEMPR0[18] ), .B(\A_DOUT_TEMPR1[18] ), .C(
        \A_DOUT_TEMPR2[18] ), .D(\A_DOUT_TEMPR3[18] ), .Y(OR4_613_Y));
    OR4 OR4_144 (.A(\A_DOUT_TEMPR79[27] ), .B(\A_DOUT_TEMPR80[27] ), 
        .C(\A_DOUT_TEMPR81[27] ), .D(\A_DOUT_TEMPR82[27] ), .Y(
        OR4_144_Y));
    OR4 OR4_2818 (.A(\B_DOUT_TEMPR52[15] ), .B(\B_DOUT_TEMPR53[15] ), 
        .C(\B_DOUT_TEMPR54[15] ), .D(\B_DOUT_TEMPR55[15] ), .Y(
        OR4_2818_Y));
    OR4 OR4_344 (.A(\B_DOUT_TEMPR79[29] ), .B(\B_DOUT_TEMPR80[29] ), 
        .C(\B_DOUT_TEMPR81[29] ), .D(\B_DOUT_TEMPR82[29] ), .Y(
        OR4_344_Y));
    OR4 OR4_826 (.A(\B_DOUT_TEMPR12[31] ), .B(\B_DOUT_TEMPR13[31] ), 
        .C(\B_DOUT_TEMPR14[31] ), .D(\B_DOUT_TEMPR15[31] ), .Y(
        OR4_826_Y));
    OR4 OR4_1474 (.A(OR4_2449_Y), .B(OR4_230_Y), .C(OR4_2319_Y), .D(
        OR4_2172_Y), .Y(OR4_1474_Y));
    OR4 OR4_1845 (.A(\B_DOUT_TEMPR40[37] ), .B(\B_DOUT_TEMPR41[37] ), 
        .C(\B_DOUT_TEMPR42[37] ), .D(\B_DOUT_TEMPR43[37] ), .Y(
        OR4_1845_Y));
    OR4 OR4_3008 (.A(\B_DOUT_TEMPR87[25] ), .B(\B_DOUT_TEMPR88[25] ), 
        .C(\B_DOUT_TEMPR89[25] ), .D(\B_DOUT_TEMPR90[25] ), .Y(
        OR4_3008_Y));
    OR4 OR4_398 (.A(\B_DOUT_TEMPR68[39] ), .B(\B_DOUT_TEMPR69[39] ), 
        .C(\B_DOUT_TEMPR70[39] ), .D(\B_DOUT_TEMPR71[39] ), .Y(
        OR4_398_Y));
    OR2 OR2_66 (.A(\A_DOUT_TEMPR72[30] ), .B(\A_DOUT_TEMPR73[30] ), .Y(
        OR2_66_Y));
    OR4 \OR4_A_DOUT[26]  (.A(OR4_1309_Y), .B(OR4_1946_Y), .C(OR4_704_Y)
        , .D(OR4_711_Y), .Y(A_DOUT[26]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%70%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R70C2 (
        .A_DOUT({nc17550, nc17551, nc17552, nc17553, nc17554, nc17555, 
        nc17556, nc17557, nc17558, nc17559, nc17560, nc17561, nc17562, 
        nc17563, nc17564, \A_DOUT_TEMPR70[14] , \A_DOUT_TEMPR70[13] , 
        \A_DOUT_TEMPR70[12] , \A_DOUT_TEMPR70[11] , 
        \A_DOUT_TEMPR70[10] }), .B_DOUT({nc17565, nc17566, nc17567, 
        nc17568, nc17569, nc17570, nc17571, nc17572, nc17573, nc17574, 
        nc17575, nc17576, nc17577, nc17578, nc17579, 
        \B_DOUT_TEMPR70[14] , \B_DOUT_TEMPR70[13] , 
        \B_DOUT_TEMPR70[12] , \B_DOUT_TEMPR70[11] , 
        \B_DOUT_TEMPR70[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[70][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_252 (.A(\B_DOUT_TEMPR103[18] ), .B(\B_DOUT_TEMPR104[18] ), 
        .C(\B_DOUT_TEMPR105[18] ), .D(\B_DOUT_TEMPR106[18] ), .Y(
        OR4_252_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%98%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R98C1 (
        .A_DOUT({nc17580, nc17581, nc17582, nc17583, nc17584, nc17585, 
        nc17586, nc17587, nc17588, nc17589, nc17590, nc17591, nc17592, 
        nc17593, nc17594, \A_DOUT_TEMPR98[9] , \A_DOUT_TEMPR98[8] , 
        \A_DOUT_TEMPR98[7] , \A_DOUT_TEMPR98[6] , \A_DOUT_TEMPR98[5] })
        , .B_DOUT({nc17595, nc17596, nc17597, nc17598, nc17599, 
        nc17600, nc17601, nc17602, nc17603, nc17604, nc17605, nc17606, 
        nc17607, nc17608, nc17609, \B_DOUT_TEMPR98[9] , 
        \B_DOUT_TEMPR98[8] , \B_DOUT_TEMPR98[7] , \B_DOUT_TEMPR98[6] , 
        \B_DOUT_TEMPR98[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[98][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%8%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R8C7 (
        .A_DOUT({nc17610, nc17611, nc17612, nc17613, nc17614, nc17615, 
        nc17616, nc17617, nc17618, nc17619, nc17620, nc17621, nc17622, 
        nc17623, nc17624, \A_DOUT_TEMPR8[39] , \A_DOUT_TEMPR8[38] , 
        \A_DOUT_TEMPR8[37] , \A_DOUT_TEMPR8[36] , \A_DOUT_TEMPR8[35] })
        , .B_DOUT({nc17625, nc17626, nc17627, nc17628, nc17629, 
        nc17630, nc17631, nc17632, nc17633, nc17634, nc17635, nc17636, 
        nc17637, nc17638, nc17639, \B_DOUT_TEMPR8[39] , 
        \B_DOUT_TEMPR8[38] , \B_DOUT_TEMPR8[37] , \B_DOUT_TEMPR8[36] , 
        \B_DOUT_TEMPR8[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_795 (.A(\B_DOUT_TEMPR32[29] ), .B(\B_DOUT_TEMPR33[29] ), 
        .C(\B_DOUT_TEMPR34[29] ), .D(\B_DOUT_TEMPR35[29] ), .Y(
        OR4_795_Y));
    OR4 OR4_320 (.A(\A_DOUT_TEMPR68[24] ), .B(\A_DOUT_TEMPR69[24] ), 
        .C(\A_DOUT_TEMPR70[24] ), .D(\A_DOUT_TEMPR71[24] ), .Y(
        OR4_320_Y));
    OR4 OR4_862 (.A(\A_DOUT_TEMPR64[25] ), .B(\A_DOUT_TEMPR65[25] ), 
        .C(\A_DOUT_TEMPR66[25] ), .D(\A_DOUT_TEMPR67[25] ), .Y(
        OR4_862_Y));
    OR4 OR4_2093 (.A(OR4_1503_Y), .B(OR4_1340_Y), .C(OR4_1283_Y), .D(
        OR4_3009_Y), .Y(OR4_2093_Y));
    OR4 OR4_2760 (.A(\B_DOUT_TEMPR16[26] ), .B(\B_DOUT_TEMPR17[26] ), 
        .C(\B_DOUT_TEMPR18[26] ), .D(\B_DOUT_TEMPR19[26] ), .Y(
        OR4_2760_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%113%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R113C5 (
        .A_DOUT({nc17640, nc17641, nc17642, nc17643, nc17644, nc17645, 
        nc17646, nc17647, nc17648, nc17649, nc17650, nc17651, nc17652, 
        nc17653, nc17654, \A_DOUT_TEMPR113[29] , \A_DOUT_TEMPR113[28] , 
        \A_DOUT_TEMPR113[27] , \A_DOUT_TEMPR113[26] , 
        \A_DOUT_TEMPR113[25] }), .B_DOUT({nc17655, nc17656, nc17657, 
        nc17658, nc17659, nc17660, nc17661, nc17662, nc17663, nc17664, 
        nc17665, nc17666, nc17667, nc17668, nc17669, 
        \B_DOUT_TEMPR113[29] , \B_DOUT_TEMPR113[28] , 
        \B_DOUT_TEMPR113[27] , \B_DOUT_TEMPR113[26] , 
        \B_DOUT_TEMPR113[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[113][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%64%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R64C4 (
        .A_DOUT({nc17670, nc17671, nc17672, nc17673, nc17674, nc17675, 
        nc17676, nc17677, nc17678, nc17679, nc17680, nc17681, nc17682, 
        nc17683, nc17684, \A_DOUT_TEMPR64[24] , \A_DOUT_TEMPR64[23] , 
        \A_DOUT_TEMPR64[22] , \A_DOUT_TEMPR64[21] , 
        \A_DOUT_TEMPR64[20] }), .B_DOUT({nc17685, nc17686, nc17687, 
        nc17688, nc17689, nc17690, nc17691, nc17692, nc17693, nc17694, 
        nc17695, nc17696, nc17697, nc17698, nc17699, 
        \B_DOUT_TEMPR64[24] , \B_DOUT_TEMPR64[23] , 
        \B_DOUT_TEMPR64[22] , \B_DOUT_TEMPR64[21] , 
        \B_DOUT_TEMPR64[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[64][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_16 (.A(\A_DOUT_TEMPR72[9] ), .B(\A_DOUT_TEMPR73[9] ), .Y(
        OR2_16_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%98%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R98C7 (
        .A_DOUT({nc17700, nc17701, nc17702, nc17703, nc17704, nc17705, 
        nc17706, nc17707, nc17708, nc17709, nc17710, nc17711, nc17712, 
        nc17713, nc17714, \A_DOUT_TEMPR98[39] , \A_DOUT_TEMPR98[38] , 
        \A_DOUT_TEMPR98[37] , \A_DOUT_TEMPR98[36] , 
        \A_DOUT_TEMPR98[35] }), .B_DOUT({nc17715, nc17716, nc17717, 
        nc17718, nc17719, nc17720, nc17721, nc17722, nc17723, nc17724, 
        nc17725, nc17726, nc17727, nc17728, nc17729, 
        \B_DOUT_TEMPR98[39] , \B_DOUT_TEMPR98[38] , 
        \B_DOUT_TEMPR98[37] , \B_DOUT_TEMPR98[36] , 
        \B_DOUT_TEMPR98[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[98][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[2]  (.A(CFG3_10_Y), .B(
        CFG3_14_Y), .Y(\BLKX2[2] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%32%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R32C7 (
        .A_DOUT({nc17730, nc17731, nc17732, nc17733, nc17734, nc17735, 
        nc17736, nc17737, nc17738, nc17739, nc17740, nc17741, nc17742, 
        nc17743, nc17744, \A_DOUT_TEMPR32[39] , \A_DOUT_TEMPR32[38] , 
        \A_DOUT_TEMPR32[37] , \A_DOUT_TEMPR32[36] , 
        \A_DOUT_TEMPR32[35] }), .B_DOUT({nc17745, nc17746, nc17747, 
        nc17748, nc17749, nc17750, nc17751, nc17752, nc17753, nc17754, 
        nc17755, nc17756, nc17757, nc17758, nc17759, 
        \B_DOUT_TEMPR32[39] , \B_DOUT_TEMPR32[38] , 
        \B_DOUT_TEMPR32[37] , \B_DOUT_TEMPR32[36] , 
        \B_DOUT_TEMPR32[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[32][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2691 (.A(\B_DOUT_TEMPR56[4] ), .B(\B_DOUT_TEMPR57[4] ), .C(
        \B_DOUT_TEMPR58[4] ), .D(\B_DOUT_TEMPR59[4] ), .Y(OR4_2691_Y));
    OR4 OR4_2284 (.A(\A_DOUT_TEMPR111[27] ), .B(\A_DOUT_TEMPR112[27] ), 
        .C(\A_DOUT_TEMPR113[27] ), .D(\A_DOUT_TEMPR114[27] ), .Y(
        OR4_2284_Y));
    OR4 OR4_1069 (.A(\B_DOUT_TEMPR115[37] ), .B(\B_DOUT_TEMPR116[37] ), 
        .C(\B_DOUT_TEMPR117[37] ), .D(\B_DOUT_TEMPR118[37] ), .Y(
        OR4_1069_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%89%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R89C7 (
        .A_DOUT({nc17760, nc17761, nc17762, nc17763, nc17764, nc17765, 
        nc17766, nc17767, nc17768, nc17769, nc17770, nc17771, nc17772, 
        nc17773, nc17774, \A_DOUT_TEMPR89[39] , \A_DOUT_TEMPR89[38] , 
        \A_DOUT_TEMPR89[37] , \A_DOUT_TEMPR89[36] , 
        \A_DOUT_TEMPR89[35] }), .B_DOUT({nc17775, nc17776, nc17777, 
        nc17778, nc17779, nc17780, nc17781, nc17782, nc17783, nc17784, 
        nc17785, nc17786, nc17787, nc17788, nc17789, 
        \B_DOUT_TEMPR89[39] , \B_DOUT_TEMPR89[38] , 
        \B_DOUT_TEMPR89[37] , \B_DOUT_TEMPR89[36] , 
        \B_DOUT_TEMPR89[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[89][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2793 (.A(\A_DOUT_TEMPR79[28] ), .B(\A_DOUT_TEMPR80[28] ), 
        .C(\A_DOUT_TEMPR81[28] ), .D(\A_DOUT_TEMPR82[28] ), .Y(
        OR4_2793_Y));
    OR4 OR4_2574 (.A(\A_DOUT_TEMPR4[10] ), .B(\A_DOUT_TEMPR5[10] ), .C(
        \A_DOUT_TEMPR6[10] ), .D(\A_DOUT_TEMPR7[10] ), .Y(OR4_2574_Y));
    OR4 OR4_1569 (.A(\A_DOUT_TEMPR115[4] ), .B(\A_DOUT_TEMPR116[4] ), 
        .C(\A_DOUT_TEMPR117[4] ), .D(\A_DOUT_TEMPR118[4] ), .Y(
        OR4_1569_Y));
    OR4 OR4_1618 (.A(\B_DOUT_TEMPR95[14] ), .B(\B_DOUT_TEMPR96[14] ), 
        .C(\B_DOUT_TEMPR97[14] ), .D(\B_DOUT_TEMPR98[14] ), .Y(
        OR4_1618_Y));
    OR4 OR4_2195 (.A(OR4_1872_Y), .B(OR4_2707_Y), .C(OR4_1737_Y), .D(
        OR4_2832_Y), .Y(OR4_2195_Y));
    OR4 OR4_6 (.A(\B_DOUT_TEMPR83[3] ), .B(\B_DOUT_TEMPR84[3] ), .C(
        \B_DOUT_TEMPR85[3] ), .D(\B_DOUT_TEMPR86[3] ), .Y(OR4_6_Y));
    OR4 OR4_998 (.A(\B_DOUT_TEMPR95[13] ), .B(\B_DOUT_TEMPR96[13] ), 
        .C(\B_DOUT_TEMPR97[13] ), .D(\B_DOUT_TEMPR98[13] ), .Y(
        OR4_998_Y));
    OR4 OR4_2083 (.A(\B_DOUT_TEMPR28[35] ), .B(\B_DOUT_TEMPR29[35] ), 
        .C(\B_DOUT_TEMPR30[35] ), .D(\B_DOUT_TEMPR31[35] ), .Y(
        OR4_2083_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%17%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R17C4 (
        .A_DOUT({nc17790, nc17791, nc17792, nc17793, nc17794, nc17795, 
        nc17796, nc17797, nc17798, nc17799, nc17800, nc17801, nc17802, 
        nc17803, nc17804, \A_DOUT_TEMPR17[24] , \A_DOUT_TEMPR17[23] , 
        \A_DOUT_TEMPR17[22] , \A_DOUT_TEMPR17[21] , 
        \A_DOUT_TEMPR17[20] }), .B_DOUT({nc17805, nc17806, nc17807, 
        nc17808, nc17809, nc17810, nc17811, nc17812, nc17813, nc17814, 
        nc17815, nc17816, nc17817, nc17818, nc17819, 
        \B_DOUT_TEMPR17[24] , \B_DOUT_TEMPR17[23] , 
        \B_DOUT_TEMPR17[22] , \B_DOUT_TEMPR17[21] , 
        \B_DOUT_TEMPR17[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2718 (.A(\A_DOUT_TEMPR8[38] ), .B(\A_DOUT_TEMPR9[38] ), .C(
        \A_DOUT_TEMPR10[38] ), .D(\A_DOUT_TEMPR11[38] ), .Y(OR4_2718_Y)
        );
    OR4 OR4_2681 (.A(OR4_564_Y), .B(OR4_2634_Y), .C(OR4_2858_Y), .D(
        OR4_2647_Y), .Y(OR4_2681_Y));
    OR4 OR4_1362 (.A(OR4_2539_Y), .B(OR4_1113_Y), .C(OR4_670_Y), .D(
        OR4_2328_Y), .Y(OR4_1362_Y));
    OR4 OR4_2304 (.A(\A_DOUT_TEMPR107[22] ), .B(\A_DOUT_TEMPR108[22] ), 
        .C(\A_DOUT_TEMPR109[22] ), .D(\A_DOUT_TEMPR110[22] ), .Y(
        OR4_2304_Y));
    OR4 OR4_1554 (.A(\B_DOUT_TEMPR48[2] ), .B(\B_DOUT_TEMPR49[2] ), .C(
        \B_DOUT_TEMPR50[2] ), .D(\B_DOUT_TEMPR51[2] ), .Y(OR4_1554_Y));
    OR4 OR4_2367 (.A(\B_DOUT_TEMPR40[22] ), .B(\B_DOUT_TEMPR41[22] ), 
        .C(\B_DOUT_TEMPR42[22] ), .D(\B_DOUT_TEMPR43[22] ), .Y(
        OR4_2367_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%100%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R100C3 (
        .A_DOUT({nc17820, nc17821, nc17822, nc17823, nc17824, nc17825, 
        nc17826, nc17827, nc17828, nc17829, nc17830, nc17831, nc17832, 
        nc17833, nc17834, \A_DOUT_TEMPR100[19] , \A_DOUT_TEMPR100[18] , 
        \A_DOUT_TEMPR100[17] , \A_DOUT_TEMPR100[16] , 
        \A_DOUT_TEMPR100[15] }), .B_DOUT({nc17835, nc17836, nc17837, 
        nc17838, nc17839, nc17840, nc17841, nc17842, nc17843, nc17844, 
        nc17845, nc17846, nc17847, nc17848, nc17849, 
        \B_DOUT_TEMPR100[19] , \B_DOUT_TEMPR100[18] , 
        \B_DOUT_TEMPR100[17] , \B_DOUT_TEMPR100[16] , 
        \B_DOUT_TEMPR100[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[100][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2262 (.A(\B_DOUT_TEMPR36[3] ), .B(\B_DOUT_TEMPR37[3] ), .C(
        \B_DOUT_TEMPR38[3] ), .D(\B_DOUT_TEMPR39[3] ), .Y(OR4_2262_Y));
    OR4 OR4_2091 (.A(\A_DOUT_TEMPR16[16] ), .B(\A_DOUT_TEMPR17[16] ), 
        .C(\A_DOUT_TEMPR18[16] ), .D(\A_DOUT_TEMPR19[16] ), .Y(
        OR4_2091_Y));
    OR4 OR4_2783 (.A(\A_DOUT_TEMPR99[18] ), .B(\A_DOUT_TEMPR100[18] ), 
        .C(\A_DOUT_TEMPR101[18] ), .D(\A_DOUT_TEMPR102[18] ), .Y(
        OR4_2783_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%103%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R103C2 (
        .A_DOUT({nc17850, nc17851, nc17852, nc17853, nc17854, nc17855, 
        nc17856, nc17857, nc17858, nc17859, nc17860, nc17861, nc17862, 
        nc17863, nc17864, \A_DOUT_TEMPR103[14] , \A_DOUT_TEMPR103[13] , 
        \A_DOUT_TEMPR103[12] , \A_DOUT_TEMPR103[11] , 
        \A_DOUT_TEMPR103[10] }), .B_DOUT({nc17865, nc17866, nc17867, 
        nc17868, nc17869, nc17870, nc17871, nc17872, nc17873, nc17874, 
        nc17875, nc17876, nc17877, nc17878, nc17879, 
        \B_DOUT_TEMPR103[14] , \B_DOUT_TEMPR103[13] , 
        \B_DOUT_TEMPR103[12] , \B_DOUT_TEMPR103[11] , 
        \B_DOUT_TEMPR103[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[103][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%27%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R27C0 (
        .A_DOUT({nc17880, nc17881, nc17882, nc17883, nc17884, nc17885, 
        nc17886, nc17887, nc17888, nc17889, nc17890, nc17891, nc17892, 
        nc17893, nc17894, \A_DOUT_TEMPR27[4] , \A_DOUT_TEMPR27[3] , 
        \A_DOUT_TEMPR27[2] , \A_DOUT_TEMPR27[1] , \A_DOUT_TEMPR27[0] })
        , .B_DOUT({nc17895, nc17896, nc17897, nc17898, nc17899, 
        nc17900, nc17901, nc17902, nc17903, nc17904, nc17905, nc17906, 
        nc17907, nc17908, nc17909, \B_DOUT_TEMPR27[4] , 
        \B_DOUT_TEMPR27[3] , \B_DOUT_TEMPR27[2] , \B_DOUT_TEMPR27[1] , 
        \B_DOUT_TEMPR27[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_186 (.A(\B_DOUT_TEMPR16[35] ), .B(\B_DOUT_TEMPR17[35] ), 
        .C(\B_DOUT_TEMPR18[35] ), .D(\B_DOUT_TEMPR19[35] ), .Y(
        OR4_186_Y));
    OR4 OR4_976 (.A(\A_DOUT_TEMPR40[33] ), .B(\A_DOUT_TEMPR41[33] ), 
        .C(\A_DOUT_TEMPR42[33] ), .D(\A_DOUT_TEMPR43[33] ), .Y(
        OR4_976_Y));
    OR4 OR4_2185 (.A(\A_DOUT_TEMPR107[17] ), .B(\A_DOUT_TEMPR108[17] ), 
        .C(\A_DOUT_TEMPR109[17] ), .D(\A_DOUT_TEMPR110[17] ), .Y(
        OR4_2185_Y));
    OR4 OR4_198 (.A(\B_DOUT_TEMPR8[11] ), .B(\B_DOUT_TEMPR9[11] ), .C(
        \B_DOUT_TEMPR10[11] ), .D(\B_DOUT_TEMPR11[11] ), .Y(OR4_198_Y));
    OR4 OR4_1280 (.A(\B_DOUT_TEMPR68[0] ), .B(\B_DOUT_TEMPR69[0] ), .C(
        \B_DOUT_TEMPR70[0] ), .D(\B_DOUT_TEMPR71[0] ), .Y(OR4_1280_Y));
    OR4 \OR4_A_DOUT[31]  (.A(OR4_1603_Y), .B(OR4_1226_Y), .C(OR4_891_Y)
        , .D(OR4_2879_Y), .Y(A_DOUT[31]));
    OR4 OR4_1274 (.A(\B_DOUT_TEMPR24[12] ), .B(\B_DOUT_TEMPR25[12] ), 
        .C(\B_DOUT_TEMPR26[12] ), .D(\B_DOUT_TEMPR27[12] ), .Y(
        OR4_1274_Y));
    OR4 OR4_2658 (.A(\A_DOUT_TEMPR115[8] ), .B(\A_DOUT_TEMPR116[8] ), 
        .C(\A_DOUT_TEMPR117[8] ), .D(\A_DOUT_TEMPR118[8] ), .Y(
        OR4_2658_Y));
    OR4 OR4_2271 (.A(\B_DOUT_TEMPR40[26] ), .B(\B_DOUT_TEMPR41[26] ), 
        .C(\B_DOUT_TEMPR42[26] ), .D(\B_DOUT_TEMPR43[26] ), .Y(
        OR4_2271_Y));
    OR4 OR4_846 (.A(\B_DOUT_TEMPR95[21] ), .B(\B_DOUT_TEMPR96[21] ), 
        .C(\B_DOUT_TEMPR97[21] ), .D(\B_DOUT_TEMPR98[21] ), .Y(
        OR4_846_Y));
    OR4 OR4_813 (.A(\A_DOUT_TEMPR60[3] ), .B(\A_DOUT_TEMPR61[3] ), .C(
        \A_DOUT_TEMPR62[3] ), .D(\A_DOUT_TEMPR63[3] ), .Y(OR4_813_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%13%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R13C6 (
        .A_DOUT({nc17910, nc17911, nc17912, nc17913, nc17914, nc17915, 
        nc17916, nc17917, nc17918, nc17919, nc17920, nc17921, nc17922, 
        nc17923, nc17924, \A_DOUT_TEMPR13[34] , \A_DOUT_TEMPR13[33] , 
        \A_DOUT_TEMPR13[32] , \A_DOUT_TEMPR13[31] , 
        \A_DOUT_TEMPR13[30] }), .B_DOUT({nc17925, nc17926, nc17927, 
        nc17928, nc17929, nc17930, nc17931, nc17932, nc17933, nc17934, 
        nc17935, nc17936, nc17937, nc17938, nc17939, 
        \B_DOUT_TEMPR13[34] , \B_DOUT_TEMPR13[33] , 
        \B_DOUT_TEMPR13[32] , \B_DOUT_TEMPR13[31] , 
        \B_DOUT_TEMPR13[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_399 (.A(\B_DOUT_TEMPR0[22] ), .B(\B_DOUT_TEMPR1[22] ), .C(
        \B_DOUT_TEMPR2[22] ), .D(\B_DOUT_TEMPR3[22] ), .Y(OR4_399_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%3%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R3C7 (
        .A_DOUT({nc17940, nc17941, nc17942, nc17943, nc17944, nc17945, 
        nc17946, nc17947, nc17948, nc17949, nc17950, nc17951, nc17952, 
        nc17953, nc17954, \A_DOUT_TEMPR3[39] , \A_DOUT_TEMPR3[38] , 
        \A_DOUT_TEMPR3[37] , \A_DOUT_TEMPR3[36] , \A_DOUT_TEMPR3[35] })
        , .B_DOUT({nc17955, nc17956, nc17957, nc17958, nc17959, 
        nc17960, nc17961, nc17962, nc17963, nc17964, nc17965, nc17966, 
        nc17967, nc17968, nc17969, \B_DOUT_TEMPR3[39] , 
        \B_DOUT_TEMPR3[38] , \B_DOUT_TEMPR3[37] , \B_DOUT_TEMPR3[36] , 
        \B_DOUT_TEMPR3[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%91%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R91C1 (
        .A_DOUT({nc17970, nc17971, nc17972, nc17973, nc17974, nc17975, 
        nc17976, nc17977, nc17978, nc17979, nc17980, nc17981, nc17982, 
        nc17983, nc17984, \A_DOUT_TEMPR91[9] , \A_DOUT_TEMPR91[8] , 
        \A_DOUT_TEMPR91[7] , \A_DOUT_TEMPR91[6] , \A_DOUT_TEMPR91[5] })
        , .B_DOUT({nc17985, nc17986, nc17987, nc17988, nc17989, 
        nc17990, nc17991, nc17992, nc17993, nc17994, nc17995, nc17996, 
        nc17997, nc17998, nc17999, \B_DOUT_TEMPR91[9] , 
        \B_DOUT_TEMPR91[8] , \B_DOUT_TEMPR91[7] , \B_DOUT_TEMPR91[6] , 
        \B_DOUT_TEMPR91[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[91][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2640 (.A(\A_DOUT_TEMPR87[0] ), .B(\A_DOUT_TEMPR88[0] ), .C(
        \A_DOUT_TEMPR89[0] ), .D(\A_DOUT_TEMPR90[0] ), .Y(OR4_2640_Y));
    CFG3 #( .INIT(8'h1) )  CFG3_17 (.A(A_ADDR[16]), .B(A_ADDR[15]), .C(
        A_ADDR[14]), .Y(CFG3_17_Y));
    OR4 OR4_340 (.A(\B_DOUT_TEMPR0[36] ), .B(\B_DOUT_TEMPR1[36] ), .C(
        \B_DOUT_TEMPR2[36] ), .D(\B_DOUT_TEMPR3[36] ), .Y(OR4_340_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%3%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R3C0 (
        .A_DOUT({nc18000, nc18001, nc18002, nc18003, nc18004, nc18005, 
        nc18006, nc18007, nc18008, nc18009, nc18010, nc18011, nc18012, 
        nc18013, nc18014, \A_DOUT_TEMPR3[4] , \A_DOUT_TEMPR3[3] , 
        \A_DOUT_TEMPR3[2] , \A_DOUT_TEMPR3[1] , \A_DOUT_TEMPR3[0] }), 
        .B_DOUT({nc18015, nc18016, nc18017, nc18018, nc18019, nc18020, 
        nc18021, nc18022, nc18023, nc18024, nc18025, nc18026, nc18027, 
        nc18028, nc18029, \B_DOUT_TEMPR3[4] , \B_DOUT_TEMPR3[3] , 
        \B_DOUT_TEMPR3[2] , \B_DOUT_TEMPR3[1] , \B_DOUT_TEMPR3[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[3][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[0] , A_ADDR[13], A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[0] , B_ADDR[13], B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%48%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R48C0 (
        .A_DOUT({nc18030, nc18031, nc18032, nc18033, nc18034, nc18035, 
        nc18036, nc18037, nc18038, nc18039, nc18040, nc18041, nc18042, 
        nc18043, nc18044, \A_DOUT_TEMPR48[4] , \A_DOUT_TEMPR48[3] , 
        \A_DOUT_TEMPR48[2] , \A_DOUT_TEMPR48[1] , \A_DOUT_TEMPR48[0] })
        , .B_DOUT({nc18045, nc18046, nc18047, nc18048, nc18049, 
        nc18050, nc18051, nc18052, nc18053, nc18054, nc18055, nc18056, 
        nc18057, nc18058, nc18059, \B_DOUT_TEMPR48[4] , 
        \B_DOUT_TEMPR48[3] , \B_DOUT_TEMPR48[2] , \B_DOUT_TEMPR48[1] , 
        \B_DOUT_TEMPR48[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[48][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2464 (.A(\A_DOUT_TEMPR99[9] ), .B(\A_DOUT_TEMPR100[9] ), 
        .C(\A_DOUT_TEMPR101[9] ), .D(\A_DOUT_TEMPR102[9] ), .Y(
        OR4_2464_Y));
    OR4 OR4_2048 (.A(\A_DOUT_TEMPR8[22] ), .B(\A_DOUT_TEMPR9[22] ), .C(
        \A_DOUT_TEMPR10[22] ), .D(\A_DOUT_TEMPR11[22] ), .Y(OR4_2048_Y)
        );
    OR4 OR4_2081 (.A(OR4_1395_Y), .B(OR4_2968_Y), .C(OR4_730_Y), .D(
        OR4_2823_Y), .Y(OR4_2081_Y));
    OR4 OR4_1073 (.A(\A_DOUT_TEMPR64[6] ), .B(\A_DOUT_TEMPR65[6] ), .C(
        \A_DOUT_TEMPR66[6] ), .D(\A_DOUT_TEMPR67[6] ), .Y(OR4_1073_Y));
    OR4 OR4_1565 (.A(\B_DOUT_TEMPR44[22] ), .B(\B_DOUT_TEMPR45[22] ), 
        .C(\B_DOUT_TEMPR46[22] ), .D(\B_DOUT_TEMPR47[22] ), .Y(
        OR4_1565_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[21]  (.A(CFG3_6_Y), .B(
        CFG3_21_Y), .Y(\BLKY2[21] ));
    OR4 OR4_1251 (.A(\B_DOUT_TEMPR36[4] ), .B(\B_DOUT_TEMPR37[4] ), .C(
        \B_DOUT_TEMPR38[4] ), .D(\B_DOUT_TEMPR39[4] ), .Y(OR4_1251_Y));
    OR4 OR4_224 (.A(\B_DOUT_TEMPR32[9] ), .B(\B_DOUT_TEMPR33[9] ), .C(
        \B_DOUT_TEMPR34[9] ), .D(\B_DOUT_TEMPR35[9] ), .Y(OR4_224_Y));
    OR4 OR4_1671 (.A(\B_DOUT_TEMPR64[1] ), .B(\B_DOUT_TEMPR65[1] ), .C(
        \B_DOUT_TEMPR66[1] ), .D(\B_DOUT_TEMPR67[1] ), .Y(OR4_1671_Y));
    OR4 OR4_1325 (.A(OR4_1222_Y), .B(OR4_2379_Y), .C(OR2_14_Y), .D(
        \B_DOUT_TEMPR74[19] ), .Y(OR4_1325_Y));
    OR4 OR4_1386 (.A(\B_DOUT_TEMPR40[33] ), .B(\B_DOUT_TEMPR41[33] ), 
        .C(\B_DOUT_TEMPR42[33] ), .D(\B_DOUT_TEMPR43[33] ), .Y(
        OR4_1386_Y));
    OR4 OR4_3027 (.A(OR4_43_Y), .B(OR4_417_Y), .C(OR4_1182_Y), .D(
        OR4_1972_Y), .Y(OR4_3027_Y));
    OR4 OR4_767 (.A(\A_DOUT_TEMPR44[19] ), .B(\A_DOUT_TEMPR45[19] ), 
        .C(\A_DOUT_TEMPR46[19] ), .D(\A_DOUT_TEMPR47[19] ), .Y(
        OR4_767_Y));
    OR4 OR4_583 (.A(\B_DOUT_TEMPR52[11] ), .B(\B_DOUT_TEMPR53[11] ), 
        .C(\B_DOUT_TEMPR54[11] ), .D(\B_DOUT_TEMPR55[11] ), .Y(
        OR4_583_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%74%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R74C6 (
        .A_DOUT({nc18060, nc18061, nc18062, nc18063, nc18064, nc18065, 
        nc18066, nc18067, nc18068, nc18069, nc18070, nc18071, nc18072, 
        nc18073, nc18074, \A_DOUT_TEMPR74[34] , \A_DOUT_TEMPR74[33] , 
        \A_DOUT_TEMPR74[32] , \A_DOUT_TEMPR74[31] , 
        \A_DOUT_TEMPR74[30] }), .B_DOUT({nc18075, nc18076, nc18077, 
        nc18078, nc18079, nc18080, nc18081, nc18082, nc18083, nc18084, 
        nc18085, nc18086, nc18087, nc18088, nc18089, 
        \B_DOUT_TEMPR74[34] , \B_DOUT_TEMPR74[33] , 
        \B_DOUT_TEMPR74[32] , \B_DOUT_TEMPR74[31] , 
        \B_DOUT_TEMPR74[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[74][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1773 (.A(\B_DOUT_TEMPR36[2] ), .B(\B_DOUT_TEMPR37[2] ), .C(
        \B_DOUT_TEMPR38[2] ), .D(\B_DOUT_TEMPR39[2] ), .Y(OR4_1773_Y));
    OR4 OR4_112 (.A(\B_DOUT_TEMPR16[25] ), .B(\B_DOUT_TEMPR17[25] ), 
        .C(\B_DOUT_TEMPR18[25] ), .D(\B_DOUT_TEMPR19[25] ), .Y(
        OR4_112_Y));
    OR4 OR4_720 (.A(\B_DOUT_TEMPR44[11] ), .B(\B_DOUT_TEMPR45[11] ), 
        .C(\B_DOUT_TEMPR46[11] ), .D(\B_DOUT_TEMPR47[11] ), .Y(
        OR4_720_Y));
    OR4 OR4_363 (.A(OR4_1105_Y), .B(OR4_1464_Y), .C(OR4_2192_Y), .D(
        OR4_10_Y), .Y(OR4_363_Y));
    OR4 OR4_1175 (.A(\B_DOUT_TEMPR28[7] ), .B(\B_DOUT_TEMPR29[7] ), .C(
        \B_DOUT_TEMPR30[7] ), .D(\B_DOUT_TEMPR31[7] ), .Y(OR4_1175_Y));
    OR4 OR4_768 (.A(OR4_2929_Y), .B(OR4_1829_Y), .C(OR4_450_Y), .D(
        OR4_1439_Y), .Y(OR4_768_Y));
    OR4 OR4_292 (.A(\A_DOUT_TEMPR56[23] ), .B(\A_DOUT_TEMPR57[23] ), 
        .C(\A_DOUT_TEMPR58[23] ), .D(\A_DOUT_TEMPR59[23] ), .Y(
        OR4_292_Y));
    OR4 OR4_2220 (.A(\A_DOUT_TEMPR107[11] ), .B(\A_DOUT_TEMPR108[11] ), 
        .C(\A_DOUT_TEMPR109[11] ), .D(\A_DOUT_TEMPR110[11] ), .Y(
        OR4_2220_Y));
    OR4 OR4_4 (.A(OR4_46_Y), .B(OR4_2626_Y), .C(OR4_1793_Y), .D(
        OR4_726_Y), .Y(OR4_4_Y));
    OR4 OR4_906 (.A(OR4_1156_Y), .B(OR4_2836_Y), .C(OR4_2233_Y), .D(
        OR4_537_Y), .Y(OR4_906_Y));
    OR4 OR4_663 (.A(\A_DOUT_TEMPR44[28] ), .B(\A_DOUT_TEMPR45[28] ), 
        .C(\A_DOUT_TEMPR46[28] ), .D(\A_DOUT_TEMPR47[28] ), .Y(
        OR4_663_Y));
    OR4 OR4_915 (.A(\A_DOUT_TEMPR64[39] ), .B(\A_DOUT_TEMPR65[39] ), 
        .C(\A_DOUT_TEMPR66[39] ), .D(\A_DOUT_TEMPR67[39] ), .Y(
        OR4_915_Y));
    OR4 OR4_1398 (.A(\B_DOUT_TEMPR68[12] ), .B(\B_DOUT_TEMPR69[12] ), 
        .C(\B_DOUT_TEMPR70[12] ), .D(\B_DOUT_TEMPR71[12] ), .Y(
        OR4_1398_Y));
    OR4 OR4_415 (.A(\B_DOUT_TEMPR40[4] ), .B(\B_DOUT_TEMPR41[4] ), .C(
        \B_DOUT_TEMPR42[4] ), .D(\B_DOUT_TEMPR43[4] ), .Y(OR4_415_Y));
    OR4 OR4_2731 (.A(\B_DOUT_TEMPR107[32] ), .B(\B_DOUT_TEMPR108[32] ), 
        .C(\B_DOUT_TEMPR109[32] ), .D(\B_DOUT_TEMPR110[32] ), .Y(
        OR4_2731_Y));
    OR4 OR4_1102 (.A(\A_DOUT_TEMPR36[8] ), .B(\A_DOUT_TEMPR37[8] ), .C(
        \A_DOUT_TEMPR38[8] ), .D(\A_DOUT_TEMPR39[8] ), .Y(OR4_1102_Y));
    OR4 OR4_1648 (.A(OR4_736_Y), .B(OR4_1072_Y), .C(OR4_681_Y), .D(
        OR4_1091_Y), .Y(OR4_1648_Y));
    OR4 OR4_1968 (.A(\B_DOUT_TEMPR103[21] ), .B(\B_DOUT_TEMPR104[21] ), 
        .C(\B_DOUT_TEMPR105[21] ), .D(\B_DOUT_TEMPR106[21] ), .Y(
        OR4_1968_Y));
    OR4 OR4_1071 (.A(\B_DOUT_TEMPR8[32] ), .B(\B_DOUT_TEMPR9[32] ), .C(
        \B_DOUT_TEMPR10[32] ), .D(\B_DOUT_TEMPR11[32] ), .Y(OR4_1071_Y)
        );
    OR4 OR4_2400 (.A(OR4_809_Y), .B(OR4_1130_Y), .C(OR4_732_Y), .D(
        OR4_1146_Y), .Y(OR4_2400_Y));
    OR4 OR4_1731 (.A(\B_DOUT_TEMPR36[22] ), .B(\B_DOUT_TEMPR37[22] ), 
        .C(\B_DOUT_TEMPR38[22] ), .D(\B_DOUT_TEMPR39[22] ), .Y(
        OR4_1731_Y));
    OR4 OR4_2144 (.A(\B_DOUT_TEMPR107[5] ), .B(\B_DOUT_TEMPR108[5] ), 
        .C(\B_DOUT_TEMPR109[5] ), .D(\B_DOUT_TEMPR110[5] ), .Y(
        OR4_2144_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%14%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R14C4 (
        .A_DOUT({nc18090, nc18091, nc18092, nc18093, nc18094, nc18095, 
        nc18096, nc18097, nc18098, nc18099, nc18100, nc18101, nc18102, 
        nc18103, nc18104, \A_DOUT_TEMPR14[24] , \A_DOUT_TEMPR14[23] , 
        \A_DOUT_TEMPR14[22] , \A_DOUT_TEMPR14[21] , 
        \A_DOUT_TEMPR14[20] }), .B_DOUT({nc18105, nc18106, nc18107, 
        nc18108, nc18109, nc18110, nc18111, nc18112, nc18113, nc18114, 
        nc18115, nc18116, nc18117, nc18118, nc18119, 
        \B_DOUT_TEMPR14[24] , \B_DOUT_TEMPR14[23] , 
        \B_DOUT_TEMPR14[22] , \B_DOUT_TEMPR14[21] , 
        \B_DOUT_TEMPR14[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%45%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R45C0 (
        .A_DOUT({nc18120, nc18121, nc18122, nc18123, nc18124, nc18125, 
        nc18126, nc18127, nc18128, nc18129, nc18130, nc18131, nc18132, 
        nc18133, nc18134, \A_DOUT_TEMPR45[4] , \A_DOUT_TEMPR45[3] , 
        \A_DOUT_TEMPR45[2] , \A_DOUT_TEMPR45[1] , \A_DOUT_TEMPR45[0] })
        , .B_DOUT({nc18135, nc18136, nc18137, nc18138, nc18139, 
        nc18140, nc18141, nc18142, nc18143, nc18144, nc18145, nc18146, 
        nc18147, nc18148, nc18149, \B_DOUT_TEMPR45[4] , 
        \B_DOUT_TEMPR45[3] , \B_DOUT_TEMPR45[2] , \B_DOUT_TEMPR45[1] , 
        \B_DOUT_TEMPR45[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%62%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R62C7 (
        .A_DOUT({nc18150, nc18151, nc18152, nc18153, nc18154, nc18155, 
        nc18156, nc18157, nc18158, nc18159, nc18160, nc18161, nc18162, 
        nc18163, nc18164, \A_DOUT_TEMPR62[39] , \A_DOUT_TEMPR62[38] , 
        \A_DOUT_TEMPR62[37] , \A_DOUT_TEMPR62[36] , 
        \A_DOUT_TEMPR62[35] }), .B_DOUT({nc18165, nc18166, nc18167, 
        nc18168, nc18169, nc18170, nc18171, nc18172, nc18173, nc18174, 
        nc18175, nc18176, nc18177, nc18178, nc18179, 
        \B_DOUT_TEMPR62[39] , \B_DOUT_TEMPR62[38] , 
        \B_DOUT_TEMPR62[37] , \B_DOUT_TEMPR62[36] , 
        \B_DOUT_TEMPR62[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[62][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1819 (.A(\B_DOUT_TEMPR91[1] ), .B(\B_DOUT_TEMPR92[1] ), .C(
        \B_DOUT_TEMPR93[1] ), .D(\B_DOUT_TEMPR94[1] ), .Y(OR4_1819_Y));
    OR4 OR4_2326 (.A(OR4_2163_Y), .B(OR4_2911_Y), .C(OR4_1345_Y), .D(
        OR4_2914_Y), .Y(OR4_2326_Y));
    OR4 OR4_2264 (.A(\A_DOUT_TEMPR40[5] ), .B(\A_DOUT_TEMPR41[5] ), .C(
        \A_DOUT_TEMPR42[5] ), .D(\A_DOUT_TEMPR43[5] ), .Y(OR4_2264_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%101%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R101C5 (
        .A_DOUT({nc18180, nc18181, nc18182, nc18183, nc18184, nc18185, 
        nc18186, nc18187, nc18188, nc18189, nc18190, nc18191, nc18192, 
        nc18193, nc18194, \A_DOUT_TEMPR101[29] , \A_DOUT_TEMPR101[28] , 
        \A_DOUT_TEMPR101[27] , \A_DOUT_TEMPR101[26] , 
        \A_DOUT_TEMPR101[25] }), .B_DOUT({nc18195, nc18196, nc18197, 
        nc18198, nc18199, nc18200, nc18201, nc18202, nc18203, nc18204, 
        nc18205, nc18206, nc18207, nc18208, nc18209, 
        \B_DOUT_TEMPR101[29] , \B_DOUT_TEMPR101[28] , 
        \B_DOUT_TEMPR101[27] , \B_DOUT_TEMPR101[26] , 
        \B_DOUT_TEMPR101[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[101][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%58%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R58C1 (
        .A_DOUT({nc18210, nc18211, nc18212, nc18213, nc18214, nc18215, 
        nc18216, nc18217, nc18218, nc18219, nc18220, nc18221, nc18222, 
        nc18223, nc18224, \A_DOUT_TEMPR58[9] , \A_DOUT_TEMPR58[8] , 
        \A_DOUT_TEMPR58[7] , \A_DOUT_TEMPR58[6] , \A_DOUT_TEMPR58[5] })
        , .B_DOUT({nc18225, nc18226, nc18227, nc18228, nc18229, 
        nc18230, nc18231, nc18232, nc18233, nc18234, nc18235, nc18236, 
        nc18237, nc18238, nc18239, \B_DOUT_TEMPR58[9] , 
        \B_DOUT_TEMPR58[8] , \B_DOUT_TEMPR58[7] , \B_DOUT_TEMPR58[6] , 
        \B_DOUT_TEMPR58[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[58][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1111 (.A(\A_DOUT_TEMPR4[38] ), .B(\A_DOUT_TEMPR5[38] ), .C(
        \A_DOUT_TEMPR6[38] ), .D(\A_DOUT_TEMPR7[38] ), .Y(OR4_1111_Y));
    OR4 OR4_2205 (.A(\B_DOUT_TEMPR48[9] ), .B(\B_DOUT_TEMPR49[9] ), .C(
        \B_DOUT_TEMPR50[9] ), .D(\B_DOUT_TEMPR51[9] ), .Y(OR4_2205_Y));
    OR4 OR4_1482 (.A(\A_DOUT_TEMPR48[24] ), .B(\A_DOUT_TEMPR49[24] ), 
        .C(\A_DOUT_TEMPR50[24] ), .D(\A_DOUT_TEMPR51[24] ), .Y(
        OR4_1482_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%58%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R58C7 (
        .A_DOUT({nc18240, nc18241, nc18242, nc18243, nc18244, nc18245, 
        nc18246, nc18247, nc18248, nc18249, nc18250, nc18251, nc18252, 
        nc18253, nc18254, \A_DOUT_TEMPR58[39] , \A_DOUT_TEMPR58[38] , 
        \A_DOUT_TEMPR58[37] , \A_DOUT_TEMPR58[36] , 
        \A_DOUT_TEMPR58[35] }), .B_DOUT({nc18255, nc18256, nc18257, 
        nc18258, nc18259, nc18260, nc18261, nc18262, nc18263, nc18264, 
        nc18265, nc18266, nc18267, nc18268, nc18269, 
        \B_DOUT_TEMPR58[39] , \B_DOUT_TEMPR58[38] , 
        \B_DOUT_TEMPR58[37] , \B_DOUT_TEMPR58[36] , 
        \B_DOUT_TEMPR58[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[58][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_244 (.A(\B_DOUT_TEMPR64[5] ), .B(\B_DOUT_TEMPR65[5] ), .C(
        \B_DOUT_TEMPR66[5] ), .D(\B_DOUT_TEMPR67[5] ), .Y(OR4_244_Y));
    OR4 OR4_472 (.A(\B_DOUT_TEMPR48[28] ), .B(\B_DOUT_TEMPR49[28] ), 
        .C(\B_DOUT_TEMPR50[28] ), .D(\B_DOUT_TEMPR51[28] ), .Y(
        OR4_472_Y));
    OR4 OR4_3032 (.A(\A_DOUT_TEMPR4[29] ), .B(\A_DOUT_TEMPR5[29] ), .C(
        \A_DOUT_TEMPR6[29] ), .D(\A_DOUT_TEMPR7[29] ), .Y(OR4_3032_Y));
    OR4 OR4_1488 (.A(\A_DOUT_TEMPR111[5] ), .B(\A_DOUT_TEMPR112[5] ), 
        .C(\A_DOUT_TEMPR113[5] ), .D(\A_DOUT_TEMPR114[5] ), .Y(
        OR4_1488_Y));
    OR4 OR4_1015 (.A(\A_DOUT_TEMPR60[9] ), .B(\A_DOUT_TEMPR61[9] ), .C(
        \A_DOUT_TEMPR62[9] ), .D(\A_DOUT_TEMPR63[9] ), .Y(OR4_1015_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%102%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R102C0 (
        .A_DOUT({nc18270, nc18271, nc18272, nc18273, nc18274, nc18275, 
        nc18276, nc18277, nc18278, nc18279, nc18280, nc18281, nc18282, 
        nc18283, nc18284, \A_DOUT_TEMPR102[4] , \A_DOUT_TEMPR102[3] , 
        \A_DOUT_TEMPR102[2] , \A_DOUT_TEMPR102[1] , 
        \A_DOUT_TEMPR102[0] }), .B_DOUT({nc18285, nc18286, nc18287, 
        nc18288, nc18289, nc18290, nc18291, nc18292, nc18293, nc18294, 
        nc18295, nc18296, nc18297, nc18298, nc18299, 
        \B_DOUT_TEMPR102[4] , \B_DOUT_TEMPR102[3] , 
        \B_DOUT_TEMPR102[2] , \B_DOUT_TEMPR102[1] , 
        \B_DOUT_TEMPR102[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[102][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%114%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R114C1 (
        .A_DOUT({nc18300, nc18301, nc18302, nc18303, nc18304, nc18305, 
        nc18306, nc18307, nc18308, nc18309, nc18310, nc18311, nc18312, 
        nc18313, nc18314, \A_DOUT_TEMPR114[9] , \A_DOUT_TEMPR114[8] , 
        \A_DOUT_TEMPR114[7] , \A_DOUT_TEMPR114[6] , 
        \A_DOUT_TEMPR114[5] }), .B_DOUT({nc18315, nc18316, nc18317, 
        nc18318, nc18319, nc18320, nc18321, nc18322, nc18323, nc18324, 
        nc18325, nc18326, nc18327, nc18328, nc18329, 
        \B_DOUT_TEMPR114[9] , \B_DOUT_TEMPR114[8] , 
        \B_DOUT_TEMPR114[7] , \B_DOUT_TEMPR114[6] , 
        \B_DOUT_TEMPR114[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[114][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%29%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R29C6 (
        .A_DOUT({nc18330, nc18331, nc18332, nc18333, nc18334, nc18335, 
        nc18336, nc18337, nc18338, nc18339, nc18340, nc18341, nc18342, 
        nc18343, nc18344, \A_DOUT_TEMPR29[34] , \A_DOUT_TEMPR29[33] , 
        \A_DOUT_TEMPR29[32] , \A_DOUT_TEMPR29[31] , 
        \A_DOUT_TEMPR29[30] }), .B_DOUT({nc18345, nc18346, nc18347, 
        nc18348, nc18349, nc18350, nc18351, nc18352, nc18353, nc18354, 
        nc18355, nc18356, nc18357, nc18358, nc18359, 
        \B_DOUT_TEMPR29[34] , \B_DOUT_TEMPR29[33] , 
        \B_DOUT_TEMPR29[32] , \B_DOUT_TEMPR29[31] , 
        \B_DOUT_TEMPR29[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%2%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R2C0 (
        .A_DOUT({nc18360, nc18361, nc18362, nc18363, nc18364, nc18365, 
        nc18366, nc18367, nc18368, nc18369, nc18370, nc18371, nc18372, 
        nc18373, nc18374, \A_DOUT_TEMPR2[4] , \A_DOUT_TEMPR2[3] , 
        \A_DOUT_TEMPR2[2] , \A_DOUT_TEMPR2[1] , \A_DOUT_TEMPR2[0] }), 
        .B_DOUT({nc18375, nc18376, nc18377, nc18378, nc18379, nc18380, 
        nc18381, nc18382, nc18383, nc18384, nc18385, nc18386, nc18387, 
        nc18388, nc18389, \B_DOUT_TEMPR2[4] , \B_DOUT_TEMPR2[3] , 
        \B_DOUT_TEMPR2[2] , \B_DOUT_TEMPR2[1] , \B_DOUT_TEMPR2[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[2][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[0] , A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[0] , B_ADDR[13], \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2845 (.A(\B_DOUT_TEMPR75[30] ), .B(\B_DOUT_TEMPR76[30] ), 
        .C(\B_DOUT_TEMPR77[30] ), .D(\B_DOUT_TEMPR78[30] ), .Y(
        OR4_2845_Y));
    OR4 OR4_2063 (.A(\A_DOUT_TEMPR4[17] ), .B(\A_DOUT_TEMPR5[17] ), .C(
        \A_DOUT_TEMPR6[17] ), .D(\A_DOUT_TEMPR7[17] ), .Y(OR4_2063_Y));
    OR4 OR4_740 (.A(OR4_1908_Y), .B(OR4_1562_Y), .C(OR4_19_Y), .D(
        OR4_1564_Y), .Y(OR4_740_Y));
    OR4 OR4_2859 (.A(\B_DOUT_TEMPR24[28] ), .B(\B_DOUT_TEMPR25[28] ), 
        .C(\B_DOUT_TEMPR26[28] ), .D(\B_DOUT_TEMPR27[28] ), .Y(
        OR4_2859_Y));
    OR4 OR4_2433 (.A(\A_DOUT_TEMPR0[20] ), .B(\A_DOUT_TEMPR1[20] ), .C(
        \A_DOUT_TEMPR2[20] ), .D(\A_DOUT_TEMPR3[20] ), .Y(OR4_2433_Y));
    OR4 OR4_1167 (.A(\A_DOUT_TEMPR87[11] ), .B(\A_DOUT_TEMPR88[11] ), 
        .C(\A_DOUT_TEMPR89[11] ), .D(\A_DOUT_TEMPR90[11] ), .Y(
        OR4_1167_Y));
    OR4 OR4_2661 (.A(\B_DOUT_TEMPR4[38] ), .B(\B_DOUT_TEMPR5[38] ), .C(
        \B_DOUT_TEMPR6[38] ), .D(\B_DOUT_TEMPR7[38] ), .Y(OR4_2661_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%4%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R4C6 (
        .A_DOUT({nc18390, nc18391, nc18392, nc18393, nc18394, nc18395, 
        nc18396, nc18397, nc18398, nc18399, nc18400, nc18401, nc18402, 
        nc18403, nc18404, \A_DOUT_TEMPR4[34] , \A_DOUT_TEMPR4[33] , 
        \A_DOUT_TEMPR4[32] , \A_DOUT_TEMPR4[31] , \A_DOUT_TEMPR4[30] })
        , .B_DOUT({nc18405, nc18406, nc18407, nc18408, nc18409, 
        nc18410, nc18411, nc18412, nc18413, nc18414, nc18415, nc18416, 
        nc18417, nc18418, nc18419, \B_DOUT_TEMPR4[34] , 
        \B_DOUT_TEMPR4[33] , \B_DOUT_TEMPR4[32] , \B_DOUT_TEMPR4[31] , 
        \B_DOUT_TEMPR4[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1495 (.A(\A_DOUT_TEMPR103[22] ), .B(\A_DOUT_TEMPR104[22] ), 
        .C(\A_DOUT_TEMPR105[22] ), .D(\A_DOUT_TEMPR106[22] ), .Y(
        OR4_1495_Y));
    OR4 OR4_1664 (.A(\B_DOUT_TEMPR12[19] ), .B(\B_DOUT_TEMPR13[19] ), 
        .C(\B_DOUT_TEMPR14[19] ), .D(\B_DOUT_TEMPR15[19] ), .Y(
        OR4_1664_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%105%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R105C1 (
        .A_DOUT({nc18420, nc18421, nc18422, nc18423, nc18424, nc18425, 
        nc18426, nc18427, nc18428, nc18429, nc18430, nc18431, nc18432, 
        nc18433, nc18434, \A_DOUT_TEMPR105[9] , \A_DOUT_TEMPR105[8] , 
        \A_DOUT_TEMPR105[7] , \A_DOUT_TEMPR105[6] , 
        \A_DOUT_TEMPR105[5] }), .B_DOUT({nc18435, nc18436, nc18437, 
        nc18438, nc18439, nc18440, nc18441, nc18442, nc18443, nc18444, 
        nc18445, nc18446, nc18447, nc18448, nc18449, 
        \B_DOUT_TEMPR105[9] , \B_DOUT_TEMPR105[8] , 
        \B_DOUT_TEMPR105[7] , \B_DOUT_TEMPR105[6] , 
        \B_DOUT_TEMPR105[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[105][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1433 (.A(OR4_2788_Y), .B(OR4_2580_Y), .C(OR4_2519_Y), .D(
        OR4_1085_Y), .Y(OR4_1433_Y));
    OR4 OR4_2763 (.A(\A_DOUT_TEMPR44[10] ), .B(\A_DOUT_TEMPR45[10] ), 
        .C(\A_DOUT_TEMPR46[10] ), .D(\A_DOUT_TEMPR47[10] ), .Y(
        OR4_2763_Y));
    OR4 OR4_2119 (.A(\B_DOUT_TEMPR60[21] ), .B(\B_DOUT_TEMPR61[21] ), 
        .C(\B_DOUT_TEMPR62[21] ), .D(\B_DOUT_TEMPR63[21] ), .Y(
        OR4_2119_Y));
    OR4 OR4_2151 (.A(\A_DOUT_TEMPR60[31] ), .B(\A_DOUT_TEMPR61[31] ), 
        .C(\A_DOUT_TEMPR62[31] ), .D(\A_DOUT_TEMPR63[31] ), .Y(
        OR4_2151_Y));
    OR4 OR4_1580 (.A(\A_DOUT_TEMPR95[1] ), .B(\A_DOUT_TEMPR96[1] ), .C(
        \A_DOUT_TEMPR97[1] ), .D(\A_DOUT_TEMPR98[1] ), .Y(OR4_1580_Y));
    OR4 OR4_2165 (.A(\A_DOUT_TEMPR52[13] ), .B(\A_DOUT_TEMPR53[13] ), 
        .C(\A_DOUT_TEMPR54[13] ), .D(\A_DOUT_TEMPR55[13] ), .Y(
        OR4_2165_Y));
    OR4 OR4_1817 (.A(OR4_2354_Y), .B(OR4_515_Y), .C(OR4_1558_Y), .D(
        OR4_227_Y), .Y(OR4_1817_Y));
    OR4 OR4_863 (.A(\A_DOUT_TEMPR68[1] ), .B(\A_DOUT_TEMPR69[1] ), .C(
        \A_DOUT_TEMPR70[1] ), .D(\A_DOUT_TEMPR71[1] ), .Y(OR4_863_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%49%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R49C1 (
        .A_DOUT({nc18450, nc18451, nc18452, nc18453, nc18454, nc18455, 
        nc18456, nc18457, nc18458, nc18459, nc18460, nc18461, nc18462, 
        nc18463, nc18464, \A_DOUT_TEMPR49[9] , \A_DOUT_TEMPR49[8] , 
        \A_DOUT_TEMPR49[7] , \A_DOUT_TEMPR49[6] , \A_DOUT_TEMPR49[5] })
        , .B_DOUT({nc18465, nc18466, nc18467, nc18468, nc18469, 
        nc18470, nc18471, nc18472, nc18473, nc18474, nc18475, nc18476, 
        nc18477, nc18478, nc18479, \B_DOUT_TEMPR49[9] , 
        \B_DOUT_TEMPR49[8] , \B_DOUT_TEMPR49[7] , \B_DOUT_TEMPR49[6] , 
        \B_DOUT_TEMPR49[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2055 (.A(\B_DOUT_TEMPR48[3] ), .B(\B_DOUT_TEMPR49[3] ), .C(
        \B_DOUT_TEMPR50[3] ), .D(\B_DOUT_TEMPR51[3] ), .Y(OR4_2055_Y));
    OR4 OR4_2422 (.A(\A_DOUT_TEMPR20[10] ), .B(\A_DOUT_TEMPR21[10] ), 
        .C(\A_DOUT_TEMPR22[10] ), .D(\A_DOUT_TEMPR23[10] ), .Y(
        OR4_2422_Y));
    OR4 OR4_956 (.A(\A_DOUT_TEMPR8[13] ), .B(\A_DOUT_TEMPR9[13] ), .C(
        \A_DOUT_TEMPR10[13] ), .D(\A_DOUT_TEMPR11[13] ), .Y(OR4_956_Y));
    OR4 OR4_1796 (.A(\B_DOUT_TEMPR48[21] ), .B(\B_DOUT_TEMPR49[21] ), 
        .C(\B_DOUT_TEMPR50[21] ), .D(\B_DOUT_TEMPR51[21] ), .Y(
        OR4_1796_Y));
    OR4 OR4_2428 (.A(\A_DOUT_TEMPR60[27] ), .B(\A_DOUT_TEMPR61[27] ), 
        .C(\A_DOUT_TEMPR62[27] ), .D(\A_DOUT_TEMPR63[27] ), .Y(
        OR4_2428_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%49%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R49C2 (
        .A_DOUT({nc18480, nc18481, nc18482, nc18483, nc18484, nc18485, 
        nc18486, nc18487, nc18488, nc18489, nc18490, nc18491, nc18492, 
        nc18493, nc18494, \A_DOUT_TEMPR49[14] , \A_DOUT_TEMPR49[13] , 
        \A_DOUT_TEMPR49[12] , \A_DOUT_TEMPR49[11] , 
        \A_DOUT_TEMPR49[10] }), .B_DOUT({nc18495, nc18496, nc18497, 
        nc18498, nc18499, nc18500, nc18501, nc18502, nc18503, nc18504, 
        nc18505, nc18506, nc18507, nc18508, nc18509, 
        \B_DOUT_TEMPR49[14] , \B_DOUT_TEMPR49[13] , 
        \B_DOUT_TEMPR49[12] , \B_DOUT_TEMPR49[11] , 
        \B_DOUT_TEMPR49[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%9%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R9C7 (
        .A_DOUT({nc18510, nc18511, nc18512, nc18513, nc18514, nc18515, 
        nc18516, nc18517, nc18518, nc18519, nc18520, nc18521, nc18522, 
        nc18523, nc18524, \A_DOUT_TEMPR9[39] , \A_DOUT_TEMPR9[38] , 
        \A_DOUT_TEMPR9[37] , \A_DOUT_TEMPR9[36] , \A_DOUT_TEMPR9[35] })
        , .B_DOUT({nc18525, nc18526, nc18527, nc18528, nc18529, 
        nc18530, nc18531, nc18532, nc18533, nc18534, nc18535, nc18536, 
        nc18537, nc18538, nc18539, \B_DOUT_TEMPR9[39] , 
        \B_DOUT_TEMPR9[38] , \B_DOUT_TEMPR9[37] , \B_DOUT_TEMPR9[36] , 
        \B_DOUT_TEMPR9[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%45%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R45C1 (
        .A_DOUT({nc18540, nc18541, nc18542, nc18543, nc18544, nc18545, 
        nc18546, nc18547, nc18548, nc18549, nc18550, nc18551, nc18552, 
        nc18553, nc18554, \A_DOUT_TEMPR45[9] , \A_DOUT_TEMPR45[8] , 
        \A_DOUT_TEMPR45[7] , \A_DOUT_TEMPR45[6] , \A_DOUT_TEMPR45[5] })
        , .B_DOUT({nc18555, nc18556, nc18557, nc18558, nc18559, 
        nc18560, nc18561, nc18562, nc18563, nc18564, nc18565, nc18566, 
        nc18567, nc18568, nc18569, \B_DOUT_TEMPR45[9] , 
        \B_DOUT_TEMPR45[8] , \B_DOUT_TEMPR45[7] , \B_DOUT_TEMPR45[6] , 
        \B_DOUT_TEMPR45[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_402 (.A(\A_DOUT_TEMPR68[2] ), .B(\A_DOUT_TEMPR69[2] ), .C(
        \A_DOUT_TEMPR70[2] ), .D(\A_DOUT_TEMPR71[2] ), .Y(OR4_402_Y));
    OR4 OR4_2061 (.A(\B_DOUT_TEMPR107[27] ), .B(\B_DOUT_TEMPR108[27] ), 
        .C(\B_DOUT_TEMPR109[27] ), .D(\B_DOUT_TEMPR110[27] ), .Y(
        OR4_2061_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%27%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R27C1 (
        .A_DOUT({nc18570, nc18571, nc18572, nc18573, nc18574, nc18575, 
        nc18576, nc18577, nc18578, nc18579, nc18580, nc18581, nc18582, 
        nc18583, nc18584, \A_DOUT_TEMPR27[9] , \A_DOUT_TEMPR27[8] , 
        \A_DOUT_TEMPR27[7] , \A_DOUT_TEMPR27[6] , \A_DOUT_TEMPR27[5] })
        , .B_DOUT({nc18585, nc18586, nc18587, nc18588, nc18589, 
        nc18590, nc18591, nc18592, nc18593, nc18594, nc18595, nc18596, 
        nc18597, nc18598, nc18599, \B_DOUT_TEMPR27[9] , 
        \B_DOUT_TEMPR27[8] , \B_DOUT_TEMPR27[7] , \B_DOUT_TEMPR27[6] , 
        \B_DOUT_TEMPR27[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%38%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R38C1 (
        .A_DOUT({nc18600, nc18601, nc18602, nc18603, nc18604, nc18605, 
        nc18606, nc18607, nc18608, nc18609, nc18610, nc18611, nc18612, 
        nc18613, nc18614, \A_DOUT_TEMPR38[9] , \A_DOUT_TEMPR38[8] , 
        \A_DOUT_TEMPR38[7] , \A_DOUT_TEMPR38[6] , \A_DOUT_TEMPR38[5] })
        , .B_DOUT({nc18615, nc18616, nc18617, nc18618, nc18619, 
        nc18620, nc18621, nc18622, nc18623, nc18624, nc18625, nc18626, 
        nc18627, nc18628, nc18629, \B_DOUT_TEMPR38[9] , 
        \B_DOUT_TEMPR38[8] , \B_DOUT_TEMPR38[7] , \B_DOUT_TEMPR38[6] , 
        \B_DOUT_TEMPR38[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[38][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%51%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R51C1 (
        .A_DOUT({nc18630, nc18631, nc18632, nc18633, nc18634, nc18635, 
        nc18636, nc18637, nc18638, nc18639, nc18640, nc18641, nc18642, 
        nc18643, nc18644, \A_DOUT_TEMPR51[9] , \A_DOUT_TEMPR51[8] , 
        \A_DOUT_TEMPR51[7] , \A_DOUT_TEMPR51[6] , \A_DOUT_TEMPR51[5] })
        , .B_DOUT({nc18645, nc18646, nc18647, nc18648, nc18649, 
        nc18650, nc18651, nc18652, nc18653, nc18654, nc18655, nc18656, 
        nc18657, nc18658, nc18659, \B_DOUT_TEMPR51[9] , 
        \B_DOUT_TEMPR51[8] , \B_DOUT_TEMPR51[7] , \B_DOUT_TEMPR51[6] , 
        \B_DOUT_TEMPR51[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[51][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%38%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R38C7 (
        .A_DOUT({nc18660, nc18661, nc18662, nc18663, nc18664, nc18665, 
        nc18666, nc18667, nc18668, nc18669, nc18670, nc18671, nc18672, 
        nc18673, nc18674, \A_DOUT_TEMPR38[39] , \A_DOUT_TEMPR38[38] , 
        \A_DOUT_TEMPR38[37] , \A_DOUT_TEMPR38[36] , 
        \A_DOUT_TEMPR38[35] }), .B_DOUT({nc18675, nc18676, nc18677, 
        nc18678, nc18679, nc18680, nc18681, nc18682, nc18683, nc18684, 
        nc18685, nc18686, nc18687, nc18688, nc18689, 
        \B_DOUT_TEMPR38[39] , \B_DOUT_TEMPR38[38] , 
        \B_DOUT_TEMPR38[37] , \B_DOUT_TEMPR38[36] , 
        \B_DOUT_TEMPR38[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[38][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_162 (.A(\A_DOUT_TEMPR16[4] ), .B(\A_DOUT_TEMPR17[4] ), .C(
        \A_DOUT_TEMPR18[4] ), .D(\A_DOUT_TEMPR19[4] ), .Y(OR4_162_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%5%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R5C5 (
        .A_DOUT({nc18690, nc18691, nc18692, nc18693, nc18694, nc18695, 
        nc18696, nc18697, nc18698, nc18699, nc18700, nc18701, nc18702, 
        nc18703, nc18704, \A_DOUT_TEMPR5[29] , \A_DOUT_TEMPR5[28] , 
        \A_DOUT_TEMPR5[27] , \A_DOUT_TEMPR5[26] , \A_DOUT_TEMPR5[25] })
        , .B_DOUT({nc18705, nc18706, nc18707, nc18708, nc18709, 
        nc18710, nc18711, nc18712, nc18713, nc18714, nc18715, nc18716, 
        nc18717, nc18718, nc18719, \B_DOUT_TEMPR5[29] , 
        \B_DOUT_TEMPR5[28] , \B_DOUT_TEMPR5[27] , \B_DOUT_TEMPR5[26] , 
        \B_DOUT_TEMPR5[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2857 (.A(\B_DOUT_TEMPR75[16] ), .B(\B_DOUT_TEMPR76[16] ), 
        .C(\B_DOUT_TEMPR77[16] ), .D(\B_DOUT_TEMPR78[16] ), .Y(
        OR4_2857_Y));
    OR4 OR4_1209 (.A(\B_DOUT_TEMPR40[13] ), .B(\B_DOUT_TEMPR41[13] ), 
        .C(\B_DOUT_TEMPR42[13] ), .D(\B_DOUT_TEMPR43[13] ), .Y(
        OR4_1209_Y));
    OR4 OR4_1849 (.A(\B_DOUT_TEMPR75[10] ), .B(\B_DOUT_TEMPR76[10] ), 
        .C(\B_DOUT_TEMPR77[10] ), .D(\B_DOUT_TEMPR78[10] ), .Y(
        OR4_1849_Y));
    OR4 OR4_437 (.A(OR4_2848_Y), .B(OR4_84_Y), .C(OR4_2787_Y), .D(
        OR4_100_Y), .Y(OR4_437_Y));
    OR4 OR4_2606 (.A(\A_DOUT_TEMPR111[35] ), .B(\A_DOUT_TEMPR112[35] ), 
        .C(\A_DOUT_TEMPR113[35] ), .D(\A_DOUT_TEMPR114[35] ), .Y(
        OR4_2606_Y));
    OR4 OR4_2520 (.A(\A_DOUT_TEMPR40[17] ), .B(\A_DOUT_TEMPR41[17] ), 
        .C(\A_DOUT_TEMPR42[17] ), .D(\A_DOUT_TEMPR43[17] ), .Y(
        OR4_2520_Y));
    OR4 OR4_2100 (.A(\A_DOUT_TEMPR52[4] ), .B(\A_DOUT_TEMPR53[4] ), .C(
        \A_DOUT_TEMPR54[4] ), .D(\A_DOUT_TEMPR55[4] ), .Y(OR4_2100_Y));
    OR4 OR4_2695 (.A(\B_DOUT_TEMPR20[20] ), .B(\B_DOUT_TEMPR21[20] ), 
        .C(\B_DOUT_TEMPR22[20] ), .D(\B_DOUT_TEMPR23[20] ), .Y(
        OR4_2695_Y));
    OR4 OR4_1985 (.A(OR4_2939_Y), .B(OR4_698_Y), .C(OR2_71_Y), .D(
        \A_DOUT_TEMPR74[29] ), .Y(OR4_1985_Y));
    OR4 OR4_91 (.A(OR4_2894_Y), .B(OR4_647_Y), .C(OR2_70_Y), .D(
        \B_DOUT_TEMPR74[21] ), .Y(OR4_91_Y));
    OR4 OR4_965 (.A(\A_DOUT_TEMPR48[34] ), .B(\A_DOUT_TEMPR49[34] ), 
        .C(\A_DOUT_TEMPR50[34] ), .D(\A_DOUT_TEMPR51[34] ), .Y(
        OR4_965_Y));
    OR4 OR4_465 (.A(\B_DOUT_TEMPR28[32] ), .B(\B_DOUT_TEMPR29[32] ), 
        .C(\B_DOUT_TEMPR30[32] ), .D(\B_DOUT_TEMPR31[32] ), .Y(
        OR4_465_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%2%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R2C2 (
        .A_DOUT({nc18720, nc18721, nc18722, nc18723, nc18724, nc18725, 
        nc18726, nc18727, nc18728, nc18729, nc18730, nc18731, nc18732, 
        nc18733, nc18734, \A_DOUT_TEMPR2[14] , \A_DOUT_TEMPR2[13] , 
        \A_DOUT_TEMPR2[12] , \A_DOUT_TEMPR2[11] , \A_DOUT_TEMPR2[10] })
        , .B_DOUT({nc18735, nc18736, nc18737, nc18738, nc18739, 
        nc18740, nc18741, nc18742, nc18743, nc18744, nc18745, nc18746, 
        nc18747, nc18748, nc18749, \B_DOUT_TEMPR2[14] , 
        \B_DOUT_TEMPR2[13] , \B_DOUT_TEMPR2[12] , \B_DOUT_TEMPR2[11] , 
        \B_DOUT_TEMPR2[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[2][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1141 (.A(OR4_567_Y), .B(OR4_2540_Y), .C(OR4_1183_Y), .D(
        OR4_2136_Y), .Y(OR4_1141_Y));
    OR4 OR4_1689 (.A(OR4_113_Y), .B(OR4_1389_Y), .C(OR4_2075_Y), .D(
        OR4_2360_Y), .Y(OR4_1689_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%12%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R12C7 (
        .A_DOUT({nc18750, nc18751, nc18752, nc18753, nc18754, nc18755, 
        nc18756, nc18757, nc18758, nc18759, nc18760, nc18761, nc18762, 
        nc18763, nc18764, \A_DOUT_TEMPR12[39] , \A_DOUT_TEMPR12[38] , 
        \A_DOUT_TEMPR12[37] , \A_DOUT_TEMPR12[36] , 
        \A_DOUT_TEMPR12[35] }), .B_DOUT({nc18765, nc18766, nc18767, 
        nc18768, nc18769, nc18770, nc18771, nc18772, nc18773, nc18774, 
        nc18775, nc18776, nc18777, nc18778, nc18779, 
        \B_DOUT_TEMPR12[39] , \B_DOUT_TEMPR12[38] , 
        \B_DOUT_TEMPR12[37] , \B_DOUT_TEMPR12[36] , 
        \B_DOUT_TEMPR12[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%86%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R86C1 (
        .A_DOUT({nc18780, nc18781, nc18782, nc18783, nc18784, nc18785, 
        nc18786, nc18787, nc18788, nc18789, nc18790, nc18791, nc18792, 
        nc18793, nc18794, \A_DOUT_TEMPR86[9] , \A_DOUT_TEMPR86[8] , 
        \A_DOUT_TEMPR86[7] , \A_DOUT_TEMPR86[6] , \A_DOUT_TEMPR86[5] })
        , .B_DOUT({nc18795, nc18796, nc18797, nc18798, nc18799, 
        nc18800, nc18801, nc18802, nc18803, nc18804, nc18805, nc18806, 
        nc18807, nc18808, nc18809, \B_DOUT_TEMPR86[9] , 
        \B_DOUT_TEMPR86[8] , \B_DOUT_TEMPR86[7] , \B_DOUT_TEMPR86[6] , 
        \B_DOUT_TEMPR86[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[86][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1045 (.A(\B_DOUT_TEMPR48[17] ), .B(\B_DOUT_TEMPR49[17] ), 
        .C(\B_DOUT_TEMPR50[17] ), .D(\B_DOUT_TEMPR51[17] ), .Y(
        OR4_1045_Y));
    OR4 OR4_684 (.A(\B_DOUT_TEMPR64[4] ), .B(\B_DOUT_TEMPR65[4] ), .C(
        \B_DOUT_TEMPR66[4] ), .D(\B_DOUT_TEMPR67[4] ), .Y(OR4_684_Y));
    OR4 OR4_1523 (.A(\B_DOUT_TEMPR8[18] ), .B(\B_DOUT_TEMPR9[18] ), .C(
        \B_DOUT_TEMPR10[18] ), .D(\B_DOUT_TEMPR11[18] ), .Y(OR4_1523_Y)
        );
    OR4 OR4_2697 (.A(OR4_1947_Y), .B(OR4_2010_Y), .C(OR4_2724_Y), .D(
        OR4_3014_Y), .Y(OR4_2697_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%78%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R78C0 (
        .A_DOUT({nc18810, nc18811, nc18812, nc18813, nc18814, nc18815, 
        nc18816, nc18817, nc18818, nc18819, nc18820, nc18821, nc18822, 
        nc18823, nc18824, \A_DOUT_TEMPR78[4] , \A_DOUT_TEMPR78[3] , 
        \A_DOUT_TEMPR78[2] , \A_DOUT_TEMPR78[1] , \A_DOUT_TEMPR78[0] })
        , .B_DOUT({nc18825, nc18826, nc18827, nc18828, nc18829, 
        nc18830, nc18831, nc18832, nc18833, nc18834, nc18835, nc18836, 
        nc18837, nc18838, nc18839, \B_DOUT_TEMPR78[4] , 
        \B_DOUT_TEMPR78[3] , \B_DOUT_TEMPR78[2] , \B_DOUT_TEMPR78[1] , 
        \B_DOUT_TEMPR78[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[78][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%6%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R6C4 (
        .A_DOUT({nc18840, nc18841, nc18842, nc18843, nc18844, nc18845, 
        nc18846, nc18847, nc18848, nc18849, nc18850, nc18851, nc18852, 
        nc18853, nc18854, \A_DOUT_TEMPR6[24] , \A_DOUT_TEMPR6[23] , 
        \A_DOUT_TEMPR6[22] , \A_DOUT_TEMPR6[21] , \A_DOUT_TEMPR6[20] })
        , .B_DOUT({nc18855, nc18856, nc18857, nc18858, nc18859, 
        nc18860, nc18861, nc18862, nc18863, nc18864, nc18865, nc18866, 
        nc18867, nc18868, nc18869, \B_DOUT_TEMPR6[24] , 
        \B_DOUT_TEMPR6[23] , \B_DOUT_TEMPR6[22] , \B_DOUT_TEMPR6[21] , 
        \B_DOUT_TEMPR6[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2685 (.A(\B_DOUT_TEMPR103[6] ), .B(\B_DOUT_TEMPR104[6] ), 
        .C(\B_DOUT_TEMPR105[6] ), .D(\B_DOUT_TEMPR106[6] ), .Y(
        OR4_2685_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%47%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R47C5 (
        .A_DOUT({nc18870, nc18871, nc18872, nc18873, nc18874, nc18875, 
        nc18876, nc18877, nc18878, nc18879, nc18880, nc18881, nc18882, 
        nc18883, nc18884, \A_DOUT_TEMPR47[29] , \A_DOUT_TEMPR47[28] , 
        \A_DOUT_TEMPR47[27] , \A_DOUT_TEMPR47[26] , 
        \A_DOUT_TEMPR47[25] }), .B_DOUT({nc18885, nc18886, nc18887, 
        nc18888, nc18889, nc18890, nc18891, nc18892, nc18893, nc18894, 
        nc18895, nc18896, nc18897, nc18898, nc18899, 
        \B_DOUT_TEMPR47[29] , \B_DOUT_TEMPR47[28] , 
        \B_DOUT_TEMPR47[27] , \B_DOUT_TEMPR47[26] , 
        \B_DOUT_TEMPR47[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2236 (.A(\B_DOUT_TEMPR79[0] ), .B(\B_DOUT_TEMPR80[0] ), .C(
        \B_DOUT_TEMPR81[0] ), .D(\B_DOUT_TEMPR82[0] ), .Y(OR4_2236_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%93%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R93C2 (
        .A_DOUT({nc18900, nc18901, nc18902, nc18903, nc18904, nc18905, 
        nc18906, nc18907, nc18908, nc18909, nc18910, nc18911, nc18912, 
        nc18913, nc18914, \A_DOUT_TEMPR93[14] , \A_DOUT_TEMPR93[13] , 
        \A_DOUT_TEMPR93[12] , \A_DOUT_TEMPR93[11] , 
        \A_DOUT_TEMPR93[10] }), .B_DOUT({nc18915, nc18916, nc18917, 
        nc18918, nc18919, nc18920, nc18921, nc18922, nc18923, nc18924, 
        nc18925, nc18926, nc18927, nc18928, nc18929, 
        \B_DOUT_TEMPR93[14] , \B_DOUT_TEMPR93[13] , 
        \B_DOUT_TEMPR93[12] , \B_DOUT_TEMPR93[11] , 
        \B_DOUT_TEMPR93[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[93][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%115%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R115C3 (
        .A_DOUT({nc18930, nc18931, nc18932, nc18933, nc18934, nc18935, 
        nc18936, nc18937, nc18938, nc18939, nc18940, nc18941, nc18942, 
        nc18943, nc18944, \A_DOUT_TEMPR115[19] , \A_DOUT_TEMPR115[18] , 
        \A_DOUT_TEMPR115[17] , \A_DOUT_TEMPR115[16] , 
        \A_DOUT_TEMPR115[15] }), .B_DOUT({nc18945, nc18946, nc18947, 
        nc18948, nc18949, nc18950, nc18951, nc18952, nc18953, nc18954, 
        nc18955, nc18956, nc18957, nc18958, nc18959, 
        \B_DOUT_TEMPR115[19] , \B_DOUT_TEMPR115[18] , 
        \B_DOUT_TEMPR115[17] , \B_DOUT_TEMPR115[16] , 
        \B_DOUT_TEMPR115[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[115][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1123 (.A(\A_DOUT_TEMPR16[23] ), .B(\A_DOUT_TEMPR17[23] ), 
        .C(\A_DOUT_TEMPR18[23] ), .D(\A_DOUT_TEMPR19[23] ), .Y(
        OR4_1123_Y));
    OR4 OR4_2812 (.A(\B_DOUT_TEMPR115[39] ), .B(\B_DOUT_TEMPR116[39] ), 
        .C(\B_DOUT_TEMPR117[39] ), .D(\B_DOUT_TEMPR118[39] ), .Y(
        OR4_2812_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[18]  (.A(CFG3_22_Y), .B(
        CFG3_21_Y), .Y(\BLKY2[18] ));
    OR4 OR4_1660 (.A(\B_DOUT_TEMPR16[34] ), .B(\B_DOUT_TEMPR17[34] ), 
        .C(\B_DOUT_TEMPR18[34] ), .D(\B_DOUT_TEMPR19[34] ), .Y(
        OR4_1660_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%86%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R86C2 (
        .A_DOUT({nc18960, nc18961, nc18962, nc18963, nc18964, nc18965, 
        nc18966, nc18967, nc18968, nc18969, nc18970, nc18971, nc18972, 
        nc18973, nc18974, \A_DOUT_TEMPR86[14] , \A_DOUT_TEMPR86[13] , 
        \A_DOUT_TEMPR86[12] , \A_DOUT_TEMPR86[11] , 
        \A_DOUT_TEMPR86[10] }), .B_DOUT({nc18975, nc18976, nc18977, 
        nc18978, nc18979, nc18980, nc18981, nc18982, nc18983, nc18984, 
        nc18985, nc18986, nc18987, nc18988, nc18989, 
        \B_DOUT_TEMPR86[14] , \B_DOUT_TEMPR86[13] , 
        \B_DOUT_TEMPR86[12] , \B_DOUT_TEMPR86[11] , 
        \B_DOUT_TEMPR86[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[86][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1236 (.A(\A_DOUT_TEMPR75[7] ), .B(\A_DOUT_TEMPR76[7] ), .C(
        \A_DOUT_TEMPR77[7] ), .D(\A_DOUT_TEMPR78[7] ), .Y(OR4_1236_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%31%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R31C1 (
        .A_DOUT({nc18990, nc18991, nc18992, nc18993, nc18994, nc18995, 
        nc18996, nc18997, nc18998, nc18999, nc19000, nc19001, nc19002, 
        nc19003, nc19004, \A_DOUT_TEMPR31[9] , \A_DOUT_TEMPR31[8] , 
        \A_DOUT_TEMPR31[7] , \A_DOUT_TEMPR31[6] , \A_DOUT_TEMPR31[5] })
        , .B_DOUT({nc19005, nc19006, nc19007, nc19008, nc19009, 
        nc19010, nc19011, nc19012, nc19013, nc19014, nc19015, nc19016, 
        nc19017, nc19018, nc19019, \B_DOUT_TEMPR31[9] , 
        \B_DOUT_TEMPR31[8] , \B_DOUT_TEMPR31[7] , \B_DOUT_TEMPR31[6] , 
        \B_DOUT_TEMPR31[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%80%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R80C6 (
        .A_DOUT({nc19020, nc19021, nc19022, nc19023, nc19024, nc19025, 
        nc19026, nc19027, nc19028, nc19029, nc19030, nc19031, nc19032, 
        nc19033, nc19034, \A_DOUT_TEMPR80[34] , \A_DOUT_TEMPR80[33] , 
        \A_DOUT_TEMPR80[32] , \A_DOUT_TEMPR80[31] , 
        \A_DOUT_TEMPR80[30] }), .B_DOUT({nc19035, nc19036, nc19037, 
        nc19038, nc19039, nc19040, nc19041, nc19042, nc19043, nc19044, 
        nc19045, nc19046, nc19047, nc19048, nc19049, 
        \B_DOUT_TEMPR80[34] , \B_DOUT_TEMPR80[33] , 
        \B_DOUT_TEMPR80[32] , \B_DOUT_TEMPR80[31] , 
        \B_DOUT_TEMPR80[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[80][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1022 (.A(OR4_2478_Y), .B(OR4_640_Y), .C(OR2_41_Y), .D(
        \A_DOUT_TEMPR74[15] ), .Y(OR4_1022_Y));
    OR4 OR4_1068 (.A(OR4_1745_Y), .B(OR4_464_Y), .C(OR4_1945_Y), .D(
        OR4_467_Y), .Y(OR4_1068_Y));
    OR4 \OR4_A_DOUT[24]  (.A(OR4_1535_Y), .B(OR4_136_Y), .C(OR4_314_Y), 
        .D(OR4_1572_Y), .Y(A_DOUT[24]));
    OR4 OR4_2925 (.A(\A_DOUT_TEMPR16[7] ), .B(\A_DOUT_TEMPR17[7] ), .C(
        \A_DOUT_TEMPR18[7] ), .D(\A_DOUT_TEMPR19[7] ), .Y(OR4_2925_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%80%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R80C5 (
        .A_DOUT({nc19050, nc19051, nc19052, nc19053, nc19054, nc19055, 
        nc19056, nc19057, nc19058, nc19059, nc19060, nc19061, nc19062, 
        nc19063, nc19064, \A_DOUT_TEMPR80[29] , \A_DOUT_TEMPR80[28] , 
        \A_DOUT_TEMPR80[27] , \A_DOUT_TEMPR80[26] , 
        \A_DOUT_TEMPR80[25] }), .B_DOUT({nc19065, nc19066, nc19067, 
        nc19068, nc19069, nc19070, nc19071, nc19072, nc19073, nc19074, 
        nc19075, nc19076, nc19077, nc19078, nc19079, 
        \B_DOUT_TEMPR80[29] , \B_DOUT_TEMPR80[28] , 
        \B_DOUT_TEMPR80[27] , \B_DOUT_TEMPR80[26] , 
        \B_DOUT_TEMPR80[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[80][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1847 (.A(\B_DOUT_TEMPR107[0] ), .B(\B_DOUT_TEMPR108[0] ), 
        .C(\B_DOUT_TEMPR109[0] ), .D(\B_DOUT_TEMPR110[0] ), .Y(
        OR4_1847_Y));
    OR4 OR4_126 (.A(\A_DOUT_TEMPR91[10] ), .B(\A_DOUT_TEMPR92[10] ), 
        .C(\A_DOUT_TEMPR93[10] ), .D(\A_DOUT_TEMPR94[10] ), .Y(
        OR4_126_Y));
    OR4 OR4_2648 (.A(\B_DOUT_TEMPR91[3] ), .B(\B_DOUT_TEMPR92[3] ), .C(
        \B_DOUT_TEMPR93[3] ), .D(\B_DOUT_TEMPR94[3] ), .Y(OR4_2648_Y));
    OR4 OR4_2687 (.A(\B_DOUT_TEMPR68[23] ), .B(\B_DOUT_TEMPR69[23] ), 
        .C(\B_DOUT_TEMPR70[23] ), .D(\B_DOUT_TEMPR71[23] ), .Y(
        OR4_2687_Y));
    OR4 OR4_2629 (.A(\B_DOUT_TEMPR60[13] ), .B(\B_DOUT_TEMPR61[13] ), 
        .C(\B_DOUT_TEMPR62[13] ), .D(\B_DOUT_TEMPR63[13] ), .Y(
        OR4_2629_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%5%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R5C2 (
        .A_DOUT({nc19080, nc19081, nc19082, nc19083, nc19084, nc19085, 
        nc19086, nc19087, nc19088, nc19089, nc19090, nc19091, nc19092, 
        nc19093, nc19094, \A_DOUT_TEMPR5[14] , \A_DOUT_TEMPR5[13] , 
        \A_DOUT_TEMPR5[12] , \A_DOUT_TEMPR5[11] , \A_DOUT_TEMPR5[10] })
        , .B_DOUT({nc19095, nc19096, nc19097, nc19098, nc19099, 
        nc19100, nc19101, nc19102, nc19103, nc19104, nc19105, nc19106, 
        nc19107, nc19108, nc19109, \B_DOUT_TEMPR5[14] , 
        \B_DOUT_TEMPR5[13] , \B_DOUT_TEMPR5[12] , \B_DOUT_TEMPR5[11] , 
        \B_DOUT_TEMPR5[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1597 (.A(\B_DOUT_TEMPR64[22] ), .B(\B_DOUT_TEMPR65[22] ), 
        .C(\B_DOUT_TEMPR66[22] ), .D(\B_DOUT_TEMPR67[22] ), .Y(
        OR4_1597_Y));
    OR4 OR4_452 (.A(OR4_2684_Y), .B(OR4_2984_Y), .C(OR4_2613_Y), .D(
        OR4_2998_Y), .Y(OR4_452_Y));
    OR4 OR4_619 (.A(\A_DOUT_TEMPR87[1] ), .B(\A_DOUT_TEMPR88[1] ), .C(
        \A_DOUT_TEMPR89[1] ), .D(\A_DOUT_TEMPR90[1] ), .Y(OR4_619_Y));
    OR4 OR4_2613 (.A(\A_DOUT_TEMPR56[28] ), .B(\A_DOUT_TEMPR57[28] ), 
        .C(\A_DOUT_TEMPR58[28] ), .D(\A_DOUT_TEMPR59[28] ), .Y(
        OR4_2613_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%99%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R99C4 (
        .A_DOUT({nc19110, nc19111, nc19112, nc19113, nc19114, nc19115, 
        nc19116, nc19117, nc19118, nc19119, nc19120, nc19121, nc19122, 
        nc19123, nc19124, \A_DOUT_TEMPR99[24] , \A_DOUT_TEMPR99[23] , 
        \A_DOUT_TEMPR99[22] , \A_DOUT_TEMPR99[21] , 
        \A_DOUT_TEMPR99[20] }), .B_DOUT({nc19125, nc19126, nc19127, 
        nc19128, nc19129, nc19130, nc19131, nc19132, nc19133, nc19134, 
        nc19135, nc19136, nc19137, nc19138, nc19139, 
        \B_DOUT_TEMPR99[24] , \B_DOUT_TEMPR99[23] , 
        \B_DOUT_TEMPR99[22] , \B_DOUT_TEMPR99[21] , 
        \B_DOUT_TEMPR99[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[99][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_996 (.A(\A_DOUT_TEMPR4[12] ), .B(\A_DOUT_TEMPR5[12] ), .C(
        \A_DOUT_TEMPR6[12] ), .D(\A_DOUT_TEMPR7[12] ), .Y(OR4_996_Y));
    OR4 OR4_1675 (.A(\B_DOUT_TEMPR20[19] ), .B(\B_DOUT_TEMPR21[19] ), 
        .C(\B_DOUT_TEMPR22[19] ), .D(\B_DOUT_TEMPR23[19] ), .Y(
        OR4_1675_Y));
    OR4 OR4_2919 (.A(\A_DOUT_TEMPR8[17] ), .B(\A_DOUT_TEMPR9[17] ), .C(
        \A_DOUT_TEMPR10[17] ), .D(\A_DOUT_TEMPR11[17] ), .Y(OR4_2919_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%103%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R103C7 (
        .A_DOUT({nc19140, nc19141, nc19142, nc19143, nc19144, nc19145, 
        nc19146, nc19147, nc19148, nc19149, nc19150, nc19151, nc19152, 
        nc19153, nc19154, \A_DOUT_TEMPR103[39] , \A_DOUT_TEMPR103[38] , 
        \A_DOUT_TEMPR103[37] , \A_DOUT_TEMPR103[36] , 
        \A_DOUT_TEMPR103[35] }), .B_DOUT({nc19155, nc19156, nc19157, 
        nc19158, nc19159, nc19160, nc19161, nc19162, nc19163, nc19164, 
        nc19165, nc19166, nc19167, nc19168, nc19169, 
        \B_DOUT_TEMPR103[39] , \B_DOUT_TEMPR103[38] , 
        \B_DOUT_TEMPR103[37] , \B_DOUT_TEMPR103[36] , 
        \B_DOUT_TEMPR103[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[103][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%75%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R75C0 (
        .A_DOUT({nc19170, nc19171, nc19172, nc19173, nc19174, nc19175, 
        nc19176, nc19177, nc19178, nc19179, nc19180, nc19181, nc19182, 
        nc19183, nc19184, \A_DOUT_TEMPR75[4] , \A_DOUT_TEMPR75[3] , 
        \A_DOUT_TEMPR75[2] , \A_DOUT_TEMPR75[1] , \A_DOUT_TEMPR75[0] })
        , .B_DOUT({nc19185, nc19186, nc19187, nc19188, nc19189, 
        nc19190, nc19191, nc19192, nc19193, nc19194, nc19195, nc19196, 
        nc19197, nc19198, nc19199, \B_DOUT_TEMPR75[4] , 
        \B_DOUT_TEMPR75[3] , \B_DOUT_TEMPR75[2] , \B_DOUT_TEMPR75[1] , 
        \B_DOUT_TEMPR75[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[75][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2836 (.A(\A_DOUT_TEMPR4[4] ), .B(\A_DOUT_TEMPR5[4] ), .C(
        \A_DOUT_TEMPR6[4] ), .D(\A_DOUT_TEMPR7[4] ), .Y(OR4_2836_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%45%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R45C7 (
        .A_DOUT({nc19200, nc19201, nc19202, nc19203, nc19204, nc19205, 
        nc19206, nc19207, nc19208, nc19209, nc19210, nc19211, nc19212, 
        nc19213, nc19214, \A_DOUT_TEMPR45[39] , \A_DOUT_TEMPR45[38] , 
        \A_DOUT_TEMPR45[37] , \A_DOUT_TEMPR45[36] , 
        \A_DOUT_TEMPR45[35] }), .B_DOUT({nc19215, nc19216, nc19217, 
        nc19218, nc19219, nc19220, nc19221, nc19222, nc19223, nc19224, 
        nc19225, nc19226, nc19227, nc19228, nc19229, 
        \B_DOUT_TEMPR45[39] , \B_DOUT_TEMPR45[38] , 
        \B_DOUT_TEMPR45[37] , \B_DOUT_TEMPR45[36] , 
        \B_DOUT_TEMPR45[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[45][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_877 (.A(OR4_737_Y), .B(OR4_2556_Y), .C(OR4_1028_Y), .D(
        OR4_2558_Y), .Y(OR4_877_Y));
    OR4 OR4_2903 (.A(\B_DOUT_TEMPR103[17] ), .B(\B_DOUT_TEMPR104[17] ), 
        .C(\B_DOUT_TEMPR105[17] ), .D(\B_DOUT_TEMPR106[17] ), .Y(
        OR4_2903_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%116%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R116C3 (
        .A_DOUT({nc19230, nc19231, nc19232, nc19233, nc19234, nc19235, 
        nc19236, nc19237, nc19238, nc19239, nc19240, nc19241, nc19242, 
        nc19243, nc19244, \A_DOUT_TEMPR116[19] , \A_DOUT_TEMPR116[18] , 
        \A_DOUT_TEMPR116[17] , \A_DOUT_TEMPR116[16] , 
        \A_DOUT_TEMPR116[15] }), .B_DOUT({nc19245, nc19246, nc19247, 
        nc19248, nc19249, nc19250, nc19251, nc19252, nc19253, nc19254, 
        nc19255, nc19256, nc19257, nc19258, nc19259, 
        \B_DOUT_TEMPR116[19] , \B_DOUT_TEMPR116[18] , 
        \B_DOUT_TEMPR116[17] , \B_DOUT_TEMPR116[16] , 
        \B_DOUT_TEMPR116[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[116][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[2]  (.A(CFG3_22_Y), .B(
        CFG3_16_Y), .Y(\BLKY2[2] ));
    OR4 OR4_1836 (.A(\A_DOUT_TEMPR107[6] ), .B(\A_DOUT_TEMPR108[6] ), 
        .C(\A_DOUT_TEMPR109[6] ), .D(\A_DOUT_TEMPR110[6] ), .Y(
        OR4_1836_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%104%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R104C7 (
        .A_DOUT({nc19260, nc19261, nc19262, nc19263, nc19264, nc19265, 
        nc19266, nc19267, nc19268, nc19269, nc19270, nc19271, nc19272, 
        nc19273, nc19274, \A_DOUT_TEMPR104[39] , \A_DOUT_TEMPR104[38] , 
        \A_DOUT_TEMPR104[37] , \A_DOUT_TEMPR104[36] , 
        \A_DOUT_TEMPR104[35] }), .B_DOUT({nc19275, nc19276, nc19277, 
        nc19278, nc19279, nc19280, nc19281, nc19282, nc19283, nc19284, 
        nc19285, nc19286, nc19287, nc19288, nc19289, 
        \B_DOUT_TEMPR104[39] , \B_DOUT_TEMPR104[38] , 
        \B_DOUT_TEMPR104[37] , \B_DOUT_TEMPR104[36] , 
        \B_DOUT_TEMPR104[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[104][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_913 (.A(\B_DOUT_TEMPR111[25] ), .B(\B_DOUT_TEMPR112[25] ), 
        .C(\B_DOUT_TEMPR113[25] ), .D(\B_DOUT_TEMPR114[25] ), .Y(
        OR4_913_Y));
    OR4 OR4_523 (.A(\A_DOUT_TEMPR20[32] ), .B(\A_DOUT_TEMPR21[32] ), 
        .C(\A_DOUT_TEMPR22[32] ), .D(\A_DOUT_TEMPR23[32] ), .Y(
        OR4_523_Y));
    OR4 \OR4_A_DOUT[1]  (.A(OR4_2690_Y), .B(OR4_3012_Y), .C(OR4_800_Y), 
        .D(OR4_870_Y), .Y(A_DOUT[1]));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENB[4]  (.A(B_WBYTE_EN[2]), .B(
        B_WEN), .Y(\WBYTEENB[4] ));
    OR4 OR4_2394 (.A(\A_DOUT_TEMPR28[8] ), .B(\A_DOUT_TEMPR29[8] ), .C(
        \A_DOUT_TEMPR30[8] ), .D(\A_DOUT_TEMPR31[8] ), .Y(OR4_2394_Y));
    OR4 OR4_1164 (.A(\A_DOUT_TEMPR79[15] ), .B(\A_DOUT_TEMPR80[15] ), 
        .C(\A_DOUT_TEMPR81[15] ), .D(\A_DOUT_TEMPR82[15] ), .Y(
        OR4_1164_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%68%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R68C1 (
        .A_DOUT({nc19290, nc19291, nc19292, nc19293, nc19294, nc19295, 
        nc19296, nc19297, nc19298, nc19299, nc19300, nc19301, nc19302, 
        nc19303, nc19304, \A_DOUT_TEMPR68[9] , \A_DOUT_TEMPR68[8] , 
        \A_DOUT_TEMPR68[7] , \A_DOUT_TEMPR68[6] , \A_DOUT_TEMPR68[5] })
        , .B_DOUT({nc19305, nc19306, nc19307, nc19308, nc19309, 
        nc19310, nc19311, nc19312, nc19313, nc19314, nc19315, nc19316, 
        nc19317, nc19318, nc19319, \B_DOUT_TEMPR68[9] , 
        \B_DOUT_TEMPR68[8] , \B_DOUT_TEMPR68[7] , \B_DOUT_TEMPR68[6] , 
        \B_DOUT_TEMPR68[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[68][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1087 (.A(OR4_2640_Y), .B(OR4_937_Y), .C(OR4_558_Y), .D(
        OR4_1604_Y), .Y(OR4_1087_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%68%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R68C7 (
        .A_DOUT({nc19320, nc19321, nc19322, nc19323, nc19324, nc19325, 
        nc19326, nc19327, nc19328, nc19329, nc19330, nc19331, nc19332, 
        nc19333, nc19334, \A_DOUT_TEMPR68[39] , \A_DOUT_TEMPR68[38] , 
        \A_DOUT_TEMPR68[37] , \A_DOUT_TEMPR68[36] , 
        \A_DOUT_TEMPR68[35] }), .B_DOUT({nc19335, nc19336, nc19337, 
        nc19338, nc19339, nc19340, nc19341, nc19342, nc19343, nc19344, 
        nc19345, nc19346, nc19347, nc19348, nc19349, 
        \B_DOUT_TEMPR68[39] , \B_DOUT_TEMPR68[38] , 
        \B_DOUT_TEMPR68[37] , \B_DOUT_TEMPR68[36] , 
        \B_DOUT_TEMPR68[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[68][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[21]  (.A(OR4_2804_Y), .B(OR4_2316_Y), .C(OR4_642_Y)
        , .D(OR4_2655_Y), .Y(B_DOUT[21]));
    OR4 OR4_1677 (.A(\B_DOUT_TEMPR99[37] ), .B(\B_DOUT_TEMPR100[37] ), 
        .C(\B_DOUT_TEMPR101[37] ), .D(\B_DOUT_TEMPR102[37] ), .Y(
        OR4_1677_Y));
    OR4 OR4_1389 (.A(\A_DOUT_TEMPR36[34] ), .B(\A_DOUT_TEMPR37[34] ), 
        .C(\A_DOUT_TEMPR38[34] ), .D(\A_DOUT_TEMPR39[34] ), .Y(
        OR4_1389_Y));
    OR4 OR4_2714 (.A(\A_DOUT_TEMPR95[13] ), .B(\A_DOUT_TEMPR96[13] ), 
        .C(\A_DOUT_TEMPR97[13] ), .D(\A_DOUT_TEMPR98[13] ), .Y(
        OR4_2714_Y));
    OR4 OR4_1287 (.A(\A_DOUT_TEMPR115[26] ), .B(\A_DOUT_TEMPR116[26] ), 
        .C(\A_DOUT_TEMPR117[26] ), .D(\A_DOUT_TEMPR118[26] ), .Y(
        OR4_1287_Y));
    OR4 OR4_3005 (.A(\B_DOUT_TEMPR87[6] ), .B(\B_DOUT_TEMPR88[6] ), .C(
        \B_DOUT_TEMPR89[6] ), .D(\B_DOUT_TEMPR90[6] ), .Y(OR4_3005_Y));
    OR4 OR4_2301 (.A(\A_DOUT_TEMPR20[8] ), .B(\A_DOUT_TEMPR21[8] ), .C(
        \A_DOUT_TEMPR22[8] ), .D(\A_DOUT_TEMPR23[8] ), .Y(OR4_2301_Y));
    OR4 OR4_687 (.A(\A_DOUT_TEMPR95[33] ), .B(\A_DOUT_TEMPR96[33] ), 
        .C(\A_DOUT_TEMPR97[33] ), .D(\A_DOUT_TEMPR98[33] ), .Y(
        OR4_687_Y));
    OR4 OR4_2411 (.A(\A_DOUT_TEMPR103[27] ), .B(\A_DOUT_TEMPR104[27] ), 
        .C(\A_DOUT_TEMPR105[27] ), .D(\A_DOUT_TEMPR106[27] ), .Y(
        OR4_2411_Y));
    OR4 OR4_2801 (.A(\A_DOUT_TEMPR111[38] ), .B(\A_DOUT_TEMPR112[38] ), 
        .C(\A_DOUT_TEMPR113[38] ), .D(\A_DOUT_TEMPR114[38] ), .Y(
        OR4_2801_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%21%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R21C0 (
        .A_DOUT({nc19350, nc19351, nc19352, nc19353, nc19354, nc19355, 
        nc19356, nc19357, nc19358, nc19359, nc19360, nc19361, nc19362, 
        nc19363, nc19364, \A_DOUT_TEMPR21[4] , \A_DOUT_TEMPR21[3] , 
        \A_DOUT_TEMPR21[2] , \A_DOUT_TEMPR21[1] , \A_DOUT_TEMPR21[0] })
        , .B_DOUT({nc19365, nc19366, nc19367, nc19368, nc19369, 
        nc19370, nc19371, nc19372, nc19373, nc19374, nc19375, nc19376, 
        nc19377, nc19378, nc19379, \B_DOUT_TEMPR21[4] , 
        \B_DOUT_TEMPR21[3] , \B_DOUT_TEMPR21[2] , \B_DOUT_TEMPR21[1] , 
        \B_DOUT_TEMPR21[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2079 (.A(\B_DOUT_TEMPR107[37] ), .B(\B_DOUT_TEMPR108[37] ), 
        .C(\B_DOUT_TEMPR109[37] ), .D(\B_DOUT_TEMPR110[37] ), .Y(
        OR4_2079_Y));
    OR4 OR4_71 (.A(OR4_2776_Y), .B(OR4_1765_Y), .C(OR4_1977_Y), .D(
        OR4_1777_Y), .Y(OR4_71_Y));
    OR4 OR4_1980 (.A(\B_DOUT_TEMPR103[30] ), .B(\B_DOUT_TEMPR104[30] ), 
        .C(\B_DOUT_TEMPR105[30] ), .D(\B_DOUT_TEMPR106[30] ), .Y(
        OR4_1980_Y));
    OR4 OR4_146 (.A(\B_DOUT_TEMPR12[29] ), .B(\B_DOUT_TEMPR13[29] ), 
        .C(\B_DOUT_TEMPR14[29] ), .D(\B_DOUT_TEMPR15[29] ), .Y(
        OR4_146_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%88%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R88C5 (
        .A_DOUT({nc19380, nc19381, nc19382, nc19383, nc19384, nc19385, 
        nc19386, nc19387, nc19388, nc19389, nc19390, nc19391, nc19392, 
        nc19393, nc19394, \A_DOUT_TEMPR88[29] , \A_DOUT_TEMPR88[28] , 
        \A_DOUT_TEMPR88[27] , \A_DOUT_TEMPR88[26] , 
        \A_DOUT_TEMPR88[25] }), .B_DOUT({nc19395, nc19396, nc19397, 
        nc19398, nc19399, nc19400, nc19401, nc19402, nc19403, nc19404, 
        nc19405, nc19406, nc19407, nc19408, nc19409, 
        \B_DOUT_TEMPR88[29] , \B_DOUT_TEMPR88[28] , 
        \B_DOUT_TEMPR88[27] , \B_DOUT_TEMPR88[26] , 
        \B_DOUT_TEMPR88[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[88][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_96 (.A(\B_DOUT_TEMPR12[7] ), .B(\B_DOUT_TEMPR13[7] ), .C(
        \B_DOUT_TEMPR14[7] ), .D(\B_DOUT_TEMPR15[7] ), .Y(OR4_96_Y));
    OR4 OR4_2730 (.A(\A_DOUT_TEMPR83[15] ), .B(\A_DOUT_TEMPR84[15] ), 
        .C(\A_DOUT_TEMPR85[15] ), .D(\A_DOUT_TEMPR86[15] ), .Y(
        OR4_2730_Y));
    OR4 OR4_2384 (.A(\A_DOUT_TEMPR95[26] ), .B(\A_DOUT_TEMPR96[26] ), 
        .C(\A_DOUT_TEMPR97[26] ), .D(\A_DOUT_TEMPR98[26] ), .Y(
        OR4_2384_Y));
    OR4 OR4_2579 (.A(\A_DOUT_TEMPR111[13] ), .B(\A_DOUT_TEMPR112[13] ), 
        .C(\A_DOUT_TEMPR113[13] ), .D(\A_DOUT_TEMPR114[13] ), .Y(
        OR4_2579_Y));
    OR4 OR4_1298 (.A(\B_DOUT_TEMPR52[25] ), .B(\B_DOUT_TEMPR53[25] ), 
        .C(\B_DOUT_TEMPR54[25] ), .D(\B_DOUT_TEMPR55[25] ), .Y(
        OR4_1298_Y));
    OR4 OR4_1865 (.A(OR4_1341_Y), .B(OR4_2842_Y), .C(OR4_359_Y), .D(
        OR4_154_Y), .Y(OR4_1865_Y));
    OR4 OR4_1730 (.A(\B_DOUT_TEMPR87[13] ), .B(\B_DOUT_TEMPR88[13] ), 
        .C(\B_DOUT_TEMPR89[13] ), .D(\B_DOUT_TEMPR90[13] ), .Y(
        OR4_1730_Y));
    OR4 OR4_807 (.A(\B_DOUT_TEMPR107[15] ), .B(\B_DOUT_TEMPR108[15] ), 
        .C(\B_DOUT_TEMPR109[15] ), .D(\B_DOUT_TEMPR110[15] ), .Y(
        OR4_807_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%0%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R0C5 (
        .A_DOUT({nc19410, nc19411, nc19412, nc19413, nc19414, nc19415, 
        nc19416, nc19417, nc19418, nc19419, nc19420, nc19421, nc19422, 
        nc19423, nc19424, \A_DOUT_TEMPR0[29] , \A_DOUT_TEMPR0[28] , 
        \A_DOUT_TEMPR0[27] , \A_DOUT_TEMPR0[26] , \A_DOUT_TEMPR0[25] })
        , .B_DOUT({nc19425, nc19426, nc19427, nc19428, nc19429, 
        nc19430, nc19431, nc19432, nc19433, nc19434, nc19435, nc19436, 
        nc19437, nc19438, nc19439, \B_DOUT_TEMPR0[29] , 
        \B_DOUT_TEMPR0[28] , \B_DOUT_TEMPR0[27] , \B_DOUT_TEMPR0[26] , 
        \B_DOUT_TEMPR0[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h20) )  CFG3_1 (.A(A_ADDR[16]), .B(A_ADDR[15]), .C(
        A_ADDR[14]), .Y(CFG3_1_Y));
    OR4 \OR4_B_DOUT[22]  (.A(OR4_2699_Y), .B(OR4_429_Y), .C(OR4_2400_Y)
        , .D(OR4_2195_Y), .Y(B_DOUT[22]));
    OR4 OR4_1112 (.A(\B_DOUT_TEMPR52[23] ), .B(\B_DOUT_TEMPR53[23] ), 
        .C(\B_DOUT_TEMPR54[23] ), .D(\B_DOUT_TEMPR55[23] ), .Y(
        OR4_1112_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%79%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R79C1 (
        .A_DOUT({nc19440, nc19441, nc19442, nc19443, nc19444, nc19445, 
        nc19446, nc19447, nc19448, nc19449, nc19450, nc19451, nc19452, 
        nc19453, nc19454, \A_DOUT_TEMPR79[9] , \A_DOUT_TEMPR79[8] , 
        \A_DOUT_TEMPR79[7] , \A_DOUT_TEMPR79[6] , \A_DOUT_TEMPR79[5] })
        , .B_DOUT({nc19455, nc19456, nc19457, nc19458, nc19459, 
        nc19460, nc19461, nc19462, nc19463, nc19464, nc19465, nc19466, 
        nc19467, nc19468, nc19469, \B_DOUT_TEMPR79[9] , 
        \B_DOUT_TEMPR79[8] , \B_DOUT_TEMPR79[7] , \B_DOUT_TEMPR79[6] , 
        \B_DOUT_TEMPR79[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[79][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%107%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R107C4 (
        .A_DOUT({nc19470, nc19471, nc19472, nc19473, nc19474, nc19475, 
        nc19476, nc19477, nc19478, nc19479, nc19480, nc19481, nc19482, 
        nc19483, nc19484, \A_DOUT_TEMPR107[24] , \A_DOUT_TEMPR107[23] , 
        \A_DOUT_TEMPR107[22] , \A_DOUT_TEMPR107[21] , 
        \A_DOUT_TEMPR107[20] }), .B_DOUT({nc19485, nc19486, nc19487, 
        nc19488, nc19489, nc19490, nc19491, nc19492, nc19493, nc19494, 
        nc19495, nc19496, nc19497, nc19498, nc19499, 
        \B_DOUT_TEMPR107[24] , \B_DOUT_TEMPR107[23] , 
        \B_DOUT_TEMPR107[22] , \B_DOUT_TEMPR107[21] , 
        \B_DOUT_TEMPR107[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[107][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%111%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R111C3 (
        .A_DOUT({nc19500, nc19501, nc19502, nc19503, nc19504, nc19505, 
        nc19506, nc19507, nc19508, nc19509, nc19510, nc19511, nc19512, 
        nc19513, nc19514, \A_DOUT_TEMPR111[19] , \A_DOUT_TEMPR111[18] , 
        \A_DOUT_TEMPR111[17] , \A_DOUT_TEMPR111[16] , 
        \A_DOUT_TEMPR111[15] }), .B_DOUT({nc19515, nc19516, nc19517, 
        nc19518, nc19519, nc19520, nc19521, nc19522, nc19523, nc19524, 
        nc19525, nc19526, nc19527, nc19528, nc19529, 
        \B_DOUT_TEMPR111[19] , \B_DOUT_TEMPR111[18] , 
        \B_DOUT_TEMPR111[17] , \B_DOUT_TEMPR111[16] , 
        \B_DOUT_TEMPR111[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[111][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1059 (.A(\B_DOUT_TEMPR103[33] ), .B(\B_DOUT_TEMPR104[33] ), 
        .C(\B_DOUT_TEMPR105[33] ), .D(\B_DOUT_TEMPR106[33] ), .Y(
        OR4_1059_Y));
    OR4 OR4_2372 (.A(\A_DOUT_TEMPR83[27] ), .B(\A_DOUT_TEMPR84[27] ), 
        .C(\A_DOUT_TEMPR85[27] ), .D(\A_DOUT_TEMPR86[27] ), .Y(
        OR4_2372_Y));
    OR4 OR4_2027 (.A(OR4_780_Y), .B(OR4_2100_Y), .C(OR4_1738_Y), .D(
        OR4_2827_Y), .Y(OR4_2027_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%81%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R81C7 (
        .A_DOUT({nc19530, nc19531, nc19532, nc19533, nc19534, nc19535, 
        nc19536, nc19537, nc19538, nc19539, nc19540, nc19541, nc19542, 
        nc19543, nc19544, \A_DOUT_TEMPR81[39] , \A_DOUT_TEMPR81[38] , 
        \A_DOUT_TEMPR81[37] , \A_DOUT_TEMPR81[36] , 
        \A_DOUT_TEMPR81[35] }), .B_DOUT({nc19545, nc19546, nc19547, 
        nc19548, nc19549, nc19550, nc19551, nc19552, nc19553, nc19554, 
        nc19555, nc19556, nc19557, nc19558, nc19559, 
        \B_DOUT_TEMPR81[39] , \B_DOUT_TEMPR81[38] , 
        \B_DOUT_TEMPR81[37] , \B_DOUT_TEMPR81[36] , 
        \B_DOUT_TEMPR81[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[81][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1782 (.A(OR4_423_Y), .B(OR4_727_Y), .C(OR4_570_Y), .D(
        OR4_1109_Y), .Y(OR4_1782_Y));
    OR4 OR4_1901 (.A(\B_DOUT_TEMPR83[26] ), .B(\B_DOUT_TEMPR84[26] ), 
        .C(\B_DOUT_TEMPR85[26] ), .D(\B_DOUT_TEMPR86[26] ), .Y(
        OR4_1901_Y));
    OR4 OR4_2329 (.A(\B_DOUT_TEMPR8[39] ), .B(\B_DOUT_TEMPR9[39] ), .C(
        \B_DOUT_TEMPR10[39] ), .D(\B_DOUT_TEMPR11[39] ), .Y(OR4_2329_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%1%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R1C4 (
        .A_DOUT({nc19560, nc19561, nc19562, nc19563, nc19564, nc19565, 
        nc19566, nc19567, nc19568, nc19569, nc19570, nc19571, nc19572, 
        nc19573, nc19574, \A_DOUT_TEMPR1[24] , \A_DOUT_TEMPR1[23] , 
        \A_DOUT_TEMPR1[22] , \A_DOUT_TEMPR1[21] , \A_DOUT_TEMPR1[20] })
        , .B_DOUT({nc19575, nc19576, nc19577, nc19578, nc19579, 
        nc19580, nc19581, nc19582, nc19583, nc19584, nc19585, nc19586, 
        nc19587, nc19588, nc19589, \B_DOUT_TEMPR1[24] , 
        \B_DOUT_TEMPR1[23] , \B_DOUT_TEMPR1[22] , \B_DOUT_TEMPR1[21] , 
        \B_DOUT_TEMPR1[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1559 (.A(OR4_2205_Y), .B(OR4_166_Y), .C(OR4_880_Y), .D(
        OR4_2533_Y), .Y(OR4_1559_Y));
    OR4 OR4_2914 (.A(\A_DOUT_TEMPR83[18] ), .B(\A_DOUT_TEMPR84[18] ), 
        .C(\A_DOUT_TEMPR85[18] ), .D(\A_DOUT_TEMPR86[18] ), .Y(
        OR4_2914_Y));
    OR4 OR4_2227 (.A(\A_DOUT_TEMPR40[19] ), .B(\A_DOUT_TEMPR41[19] ), 
        .C(\A_DOUT_TEMPR42[19] ), .D(\A_DOUT_TEMPR43[19] ), .Y(
        OR4_2227_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%79%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R79C2 (
        .A_DOUT({nc19590, nc19591, nc19592, nc19593, nc19594, nc19595, 
        nc19596, nc19597, nc19598, nc19599, nc19600, nc19601, nc19602, 
        nc19603, nc19604, \A_DOUT_TEMPR79[14] , \A_DOUT_TEMPR79[13] , 
        \A_DOUT_TEMPR79[12] , \A_DOUT_TEMPR79[11] , 
        \A_DOUT_TEMPR79[10] }), .B_DOUT({nc19605, nc19606, nc19607, 
        nc19608, nc19609, nc19610, nc19611, nc19612, nc19613, nc19614, 
        nc19615, nc19616, nc19617, nc19618, nc19619, 
        \B_DOUT_TEMPR79[14] , \B_DOUT_TEMPR79[13] , 
        \B_DOUT_TEMPR79[12] , \B_DOUT_TEMPR79[11] , 
        \B_DOUT_TEMPR79[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[79][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_287 (.A(\B_DOUT_TEMPR12[9] ), .B(\B_DOUT_TEMPR13[9] ), .C(
        \B_DOUT_TEMPR14[9] ), .D(\B_DOUT_TEMPR15[9] ), .Y(OR4_287_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%75%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R75C1 (
        .A_DOUT({nc19620, nc19621, nc19622, nc19623, nc19624, nc19625, 
        nc19626, nc19627, nc19628, nc19629, nc19630, nc19631, nc19632, 
        nc19633, nc19634, \A_DOUT_TEMPR75[9] , \A_DOUT_TEMPR75[8] , 
        \A_DOUT_TEMPR75[7] , \A_DOUT_TEMPR75[6] , \A_DOUT_TEMPR75[5] })
        , .B_DOUT({nc19635, nc19636, nc19637, nc19638, nc19639, 
        nc19640, nc19641, nc19642, nc19643, nc19644, nc19645, nc19646, 
        nc19647, nc19648, nc19649, \B_DOUT_TEMPR75[9] , 
        \B_DOUT_TEMPR75[8] , \B_DOUT_TEMPR75[7] , \B_DOUT_TEMPR75[6] , 
        \B_DOUT_TEMPR75[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[75][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2665 (.A(OR4_2921_Y), .B(OR4_2225_Y), .C(OR4_1814_Y), .D(
        OR4_455_Y), .Y(OR4_2665_Y));
    OR4 OR4_2849 (.A(\A_DOUT_TEMPR107[38] ), .B(\A_DOUT_TEMPR108[38] ), 
        .C(\A_DOUT_TEMPR109[38] ), .D(\A_DOUT_TEMPR110[38] ), .Y(
        OR4_2849_Y));
    OR4 OR4_543 (.A(OR4_2850_Y), .B(OR4_141_Y), .C(OR4_784_Y), .D(
        OR4_3031_Y), .Y(OR4_543_Y));
    OR4 OR4_2916 (.A(\A_DOUT_TEMPR36[32] ), .B(\A_DOUT_TEMPR37[32] ), 
        .C(\A_DOUT_TEMPR38[32] ), .D(\A_DOUT_TEMPR39[32] ), .Y(
        OR4_2916_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%61%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R61C1 (
        .A_DOUT({nc19650, nc19651, nc19652, nc19653, nc19654, nc19655, 
        nc19656, nc19657, nc19658, nc19659, nc19660, nc19661, nc19662, 
        nc19663, nc19664, \A_DOUT_TEMPR61[9] , \A_DOUT_TEMPR61[8] , 
        \A_DOUT_TEMPR61[7] , \A_DOUT_TEMPR61[6] , \A_DOUT_TEMPR61[5] })
        , .B_DOUT({nc19665, nc19666, nc19667, nc19668, nc19669, 
        nc19670, nc19671, nc19672, nc19673, nc19674, nc19675, nc19676, 
        nc19677, nc19678, nc19679, \B_DOUT_TEMPR61[9] , 
        \B_DOUT_TEMPR61[8] , \B_DOUT_TEMPR61[7] , \B_DOUT_TEMPR61[6] , 
        \B_DOUT_TEMPR61[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[61][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%47%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R47C2 (
        .A_DOUT({nc19680, nc19681, nc19682, nc19683, nc19684, nc19685, 
        nc19686, nc19687, nc19688, nc19689, nc19690, nc19691, nc19692, 
        nc19693, nc19694, \A_DOUT_TEMPR47[14] , \A_DOUT_TEMPR47[13] , 
        \A_DOUT_TEMPR47[12] , \A_DOUT_TEMPR47[11] , 
        \A_DOUT_TEMPR47[10] }), .B_DOUT({nc19695, nc19696, nc19697, 
        nc19698, nc19699, nc19700, nc19701, nc19702, nc19703, nc19704, 
        nc19705, nc19706, nc19707, nc19708, nc19709, 
        \B_DOUT_TEMPR47[14] , \B_DOUT_TEMPR47[13] , 
        \B_DOUT_TEMPR47[12] , \B_DOUT_TEMPR47[11] , 
        \B_DOUT_TEMPR47[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2920 (.A(\A_DOUT_TEMPR68[4] ), .B(\A_DOUT_TEMPR69[4] ), .C(
        \A_DOUT_TEMPR70[4] ), .D(\A_DOUT_TEMPR71[4] ), .Y(OR4_2920_Y));
    OR4 OR4_2337 (.A(\B_DOUT_TEMPR68[36] ), .B(\B_DOUT_TEMPR69[36] ), 
        .C(\B_DOUT_TEMPR70[36] ), .D(\B_DOUT_TEMPR71[36] ), .Y(
        OR4_2337_Y));
    OR4 OR4_2232 (.A(\B_DOUT_TEMPR107[4] ), .B(\B_DOUT_TEMPR108[4] ), 
        .C(\B_DOUT_TEMPR109[4] ), .D(\B_DOUT_TEMPR110[4] ), .Y(
        OR4_2232_Y));
    OR4 OR4_471 (.A(\B_DOUT_TEMPR103[12] ), .B(\B_DOUT_TEMPR104[12] ), 
        .C(\B_DOUT_TEMPR105[12] ), .D(\B_DOUT_TEMPR106[12] ), .Y(
        OR4_471_Y));
    CFG3 #( .INIT(8'h10) )  CFG3_8 (.A(B_ADDR[16]), .B(B_ADDR[15]), .C(
        B_ADDR[14]), .Y(CFG3_8_Y));
    OR4 OR4_1374 (.A(\B_DOUT_TEMPR20[39] ), .B(\B_DOUT_TEMPR21[39] ), 
        .C(\B_DOUT_TEMPR22[39] ), .D(\B_DOUT_TEMPR23[39] ), .Y(
        OR4_1374_Y));
    OR4 OR4_492 (.A(\B_DOUT_TEMPR75[38] ), .B(\B_DOUT_TEMPR76[38] ), 
        .C(\B_DOUT_TEMPR77[38] ), .D(\B_DOUT_TEMPR78[38] ), .Y(
        OR4_492_Y));
    OR4 OR4_1352 (.A(\A_DOUT_TEMPR111[6] ), .B(\A_DOUT_TEMPR112[6] ), 
        .C(\A_DOUT_TEMPR113[6] ), .D(\A_DOUT_TEMPR114[6] ), .Y(
        OR4_1352_Y));
    OR4 OR4_2152 (.A(\A_DOUT_TEMPR60[29] ), .B(\A_DOUT_TEMPR61[29] ), 
        .C(\A_DOUT_TEMPR62[29] ), .D(\A_DOUT_TEMPR63[29] ), .Y(
        OR4_2152_Y));
    OR4 OR4_1337 (.A(OR4_1911_Y), .B(OR4_1742_Y), .C(OR4_2438_Y), .D(
        OR4_2765_Y), .Y(OR4_1337_Y));
    OR4 OR4_2490 (.A(\B_DOUT_TEMPR56[18] ), .B(\B_DOUT_TEMPR57[18] ), 
        .C(\B_DOUT_TEMPR58[18] ), .D(\B_DOUT_TEMPR59[18] ), .Y(
        OR4_2490_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%53%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R53C2 (
        .A_DOUT({nc19710, nc19711, nc19712, nc19713, nc19714, nc19715, 
        nc19716, nc19717, nc19718, nc19719, nc19720, nc19721, nc19722, 
        nc19723, nc19724, \A_DOUT_TEMPR53[14] , \A_DOUT_TEMPR53[13] , 
        \A_DOUT_TEMPR53[12] , \A_DOUT_TEMPR53[11] , 
        \A_DOUT_TEMPR53[10] }), .B_DOUT({nc19725, nc19726, nc19727, 
        nc19728, nc19729, nc19730, nc19731, nc19732, nc19733, nc19734, 
        nc19735, nc19736, nc19737, nc19738, nc19739, 
        \B_DOUT_TEMPR53[14] , \B_DOUT_TEMPR53[13] , 
        \B_DOUT_TEMPR53[12] , \B_DOUT_TEMPR53[11] , 
        \B_DOUT_TEMPR53[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[53][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1682 (.A(\B_DOUT_TEMPR20[35] ), .B(\B_DOUT_TEMPR21[35] ), 
        .C(\B_DOUT_TEMPR22[35] ), .D(\B_DOUT_TEMPR23[35] ), .Y(
        OR4_1682_Y));
    OR4 OR4_1232 (.A(\B_DOUT_TEMPR79[12] ), .B(\B_DOUT_TEMPR80[12] ), 
        .C(\B_DOUT_TEMPR81[12] ), .D(\B_DOUT_TEMPR82[12] ), .Y(
        OR4_1232_Y));
    OR4 OR4_982 (.A(OR4_653_Y), .B(OR4_2719_Y), .C(OR4_612_Y), .D(
        OR4_1816_Y), .Y(OR4_982_Y));
    OR4 OR4_1328 (.A(\A_DOUT_TEMPR8[24] ), .B(\A_DOUT_TEMPR9[24] ), .C(
        \A_DOUT_TEMPR10[24] ), .D(\A_DOUT_TEMPR11[24] ), .Y(OR4_1328_Y)
        );
    OR4 OR4_2141 (.A(\B_DOUT_TEMPR8[7] ), .B(\B_DOUT_TEMPR9[7] ), .C(
        \B_DOUT_TEMPR10[7] ), .D(\B_DOUT_TEMPR11[7] ), .Y(OR4_2141_Y));
    OR4 OR4_3024 (.A(\A_DOUT_TEMPR56[32] ), .B(\A_DOUT_TEMPR57[32] ), 
        .C(\A_DOUT_TEMPR58[32] ), .D(\A_DOUT_TEMPR59[32] ), .Y(
        OR4_3024_Y));
    OR4 OR4_185 (.A(\A_DOUT_TEMPR107[20] ), .B(\A_DOUT_TEMPR108[20] ), 
        .C(\A_DOUT_TEMPR109[20] ), .D(\A_DOUT_TEMPR110[20] ), .Y(
        OR4_185_Y));
    OR4 OR4_3026 (.A(\B_DOUT_TEMPR36[21] ), .B(\B_DOUT_TEMPR37[21] ), 
        .C(\B_DOUT_TEMPR38[21] ), .D(\B_DOUT_TEMPR39[21] ), .Y(
        OR4_3026_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%105%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R105C6 (
        .A_DOUT({nc19740, nc19741, nc19742, nc19743, nc19744, nc19745, 
        nc19746, nc19747, nc19748, nc19749, nc19750, nc19751, nc19752, 
        nc19753, nc19754, \A_DOUT_TEMPR105[34] , \A_DOUT_TEMPR105[33] , 
        \A_DOUT_TEMPR105[32] , \A_DOUT_TEMPR105[31] , 
        \A_DOUT_TEMPR105[30] }), .B_DOUT({nc19755, nc19756, nc19757, 
        nc19758, nc19759, nc19760, nc19761, nc19762, nc19763, nc19764, 
        nc19765, nc19766, nc19767, nc19768, nc19769, 
        \B_DOUT_TEMPR105[34] , \B_DOUT_TEMPR105[33] , 
        \B_DOUT_TEMPR105[32] , \B_DOUT_TEMPR105[31] , 
        \B_DOUT_TEMPR105[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[105][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2575 (.A(OR4_819_Y), .B(OR4_94_Y), .C(OR4_2736_Y), .D(
        OR4_1361_Y), .Y(OR4_2575_Y));
    OR4 OR4_2667 (.A(\B_DOUT_TEMPR111[32] ), .B(\B_DOUT_TEMPR112[32] ), 
        .C(\B_DOUT_TEMPR113[32] ), .D(\B_DOUT_TEMPR114[32] ), .Y(
        OR4_2667_Y));
    OR4 OR4_1982 (.A(\A_DOUT_TEMPR16[22] ), .B(\A_DOUT_TEMPR17[22] ), 
        .C(\A_DOUT_TEMPR18[22] ), .D(\A_DOUT_TEMPR19[22] ), .Y(
        OR4_1982_Y));
    OR4 OR4_980 (.A(\A_DOUT_TEMPR68[27] ), .B(\A_DOUT_TEMPR69[27] ), 
        .C(\A_DOUT_TEMPR70[27] ), .D(\A_DOUT_TEMPR71[27] ), .Y(
        OR4_980_Y));
    OR4 OR4_1203 (.A(\A_DOUT_TEMPR40[10] ), .B(\A_DOUT_TEMPR41[10] ), 
        .C(\A_DOUT_TEMPR42[10] ), .D(\A_DOUT_TEMPR43[10] ), .Y(
        OR4_1203_Y));
    OR4 OR4_2045 (.A(OR4_283_Y), .B(OR4_2347_Y), .C(OR4_2566_Y), .D(
        OR4_2356_Y), .Y(OR4_2045_Y));
    OR4 OR4_669 (.A(\B_DOUT_TEMPR68[31] ), .B(\B_DOUT_TEMPR69[31] ), 
        .C(\B_DOUT_TEMPR70[31] ), .D(\B_DOUT_TEMPR71[31] ), .Y(
        OR4_669_Y));
    OR4 OR4_2722 (.A(\A_DOUT_TEMPR87[24] ), .B(\A_DOUT_TEMPR88[24] ), 
        .C(\A_DOUT_TEMPR89[24] ), .D(\A_DOUT_TEMPR90[24] ), .Y(
        OR4_2722_Y));
    OR4 OR4_2434 (.A(\B_DOUT_TEMPR87[35] ), .B(\B_DOUT_TEMPR88[35] ), 
        .C(\B_DOUT_TEMPR89[35] ), .D(\B_DOUT_TEMPR90[35] ), .Y(
        OR4_2434_Y));
    OR4 OR4_2295 (.A(\A_DOUT_TEMPR87[29] ), .B(\A_DOUT_TEMPR88[29] ), 
        .C(\A_DOUT_TEMPR89[29] ), .D(\A_DOUT_TEMPR90[29] ), .Y(
        OR4_2295_Y));
    OR4 OR4_1434 (.A(\B_DOUT_TEMPR32[8] ), .B(\B_DOUT_TEMPR33[8] ), .C(
        \B_DOUT_TEMPR34[8] ), .D(\B_DOUT_TEMPR35[8] ), .Y(OR4_1434_Y));
    OR4 OR4_2480 (.A(OR4_1873_Y), .B(OR4_911_Y), .C(OR4_1119_Y), .D(
        OR4_928_Y), .Y(OR4_2480_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[25]  (.A(CFG3_5_Y), .B(
        CFG3_18_Y), .Y(\BLKX2[25] ));
    OR4 OR4_1555 (.A(\A_DOUT_TEMPR32[25] ), .B(\A_DOUT_TEMPR33[25] ), 
        .C(\A_DOUT_TEMPR34[25] ), .D(\A_DOUT_TEMPR35[25] ), .Y(
        OR4_1555_Y));
    OR4 OR4_53 (.A(\A_DOUT_TEMPR8[30] ), .B(\A_DOUT_TEMPR9[30] ), .C(
        \A_DOUT_TEMPR10[30] ), .D(\A_DOUT_TEMPR11[30] ), .Y(OR4_53_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%18%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R18C1 (
        .A_DOUT({nc19770, nc19771, nc19772, nc19773, nc19774, nc19775, 
        nc19776, nc19777, nc19778, nc19779, nc19780, nc19781, nc19782, 
        nc19783, nc19784, \A_DOUT_TEMPR18[9] , \A_DOUT_TEMPR18[8] , 
        \A_DOUT_TEMPR18[7] , \A_DOUT_TEMPR18[6] , \A_DOUT_TEMPR18[5] })
        , .B_DOUT({nc19785, nc19786, nc19787, nc19788, nc19789, 
        nc19790, nc19791, nc19792, nc19793, nc19794, nc19795, nc19796, 
        nc19797, nc19798, nc19799, \B_DOUT_TEMPR18[9] , 
        \B_DOUT_TEMPR18[8] , \B_DOUT_TEMPR18[7] , \B_DOUT_TEMPR18[6] , 
        \B_DOUT_TEMPR18[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%59%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R59C4 (
        .A_DOUT({nc19800, nc19801, nc19802, nc19803, nc19804, nc19805, 
        nc19806, nc19807, nc19808, nc19809, nc19810, nc19811, nc19812, 
        nc19813, nc19814, \A_DOUT_TEMPR59[24] , \A_DOUT_TEMPR59[23] , 
        \A_DOUT_TEMPR59[22] , \A_DOUT_TEMPR59[21] , 
        \A_DOUT_TEMPR59[20] }), .B_DOUT({nc19815, nc19816, nc19817, 
        nc19818, nc19819, nc19820, nc19821, nc19822, nc19823, nc19824, 
        nc19825, nc19826, nc19827, nc19828, nc19829, 
        \B_DOUT_TEMPR59[24] , \B_DOUT_TEMPR59[23] , 
        \B_DOUT_TEMPR59[22] , \B_DOUT_TEMPR59[21] , 
        \B_DOUT_TEMPR59[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[59][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_963 (.A(\A_DOUT_TEMPR20[25] ), .B(\A_DOUT_TEMPR21[25] ), 
        .C(\A_DOUT_TEMPR22[25] ), .D(\A_DOUT_TEMPR23[25] ), .Y(
        OR4_963_Y));
    OR4 OR4_2847 (.A(\A_DOUT_TEMPR91[36] ), .B(\A_DOUT_TEMPR92[36] ), 
        .C(\A_DOUT_TEMPR93[36] ), .D(\A_DOUT_TEMPR94[36] ), .Y(
        OR4_2847_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%77%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R77C5 (
        .A_DOUT({nc19830, nc19831, nc19832, nc19833, nc19834, nc19835, 
        nc19836, nc19837, nc19838, nc19839, nc19840, nc19841, nc19842, 
        nc19843, nc19844, \A_DOUT_TEMPR77[29] , \A_DOUT_TEMPR77[28] , 
        \A_DOUT_TEMPR77[27] , \A_DOUT_TEMPR77[26] , 
        \A_DOUT_TEMPR77[25] }), .B_DOUT({nc19845, nc19846, nc19847, 
        nc19848, nc19849, nc19850, nc19851, nc19852, nc19853, nc19854, 
        nc19855, nc19856, nc19857, nc19858, nc19859, 
        \B_DOUT_TEMPR77[29] , \B_DOUT_TEMPR77[28] , 
        \B_DOUT_TEMPR77[27] , \B_DOUT_TEMPR77[26] , 
        \B_DOUT_TEMPR77[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[77][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_416 (.A(\A_DOUT_TEMPR48[11] ), .B(\A_DOUT_TEMPR49[11] ), 
        .C(\A_DOUT_TEMPR50[11] ), .D(\A_DOUT_TEMPR51[11] ), .Y(
        OR4_416_Y));
    OR4 OR4_401 (.A(\B_DOUT_TEMPR56[28] ), .B(\B_DOUT_TEMPR57[28] ), 
        .C(\B_DOUT_TEMPR58[28] ), .D(\B_DOUT_TEMPR59[28] ), .Y(
        OR4_401_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%18%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R18C7 (
        .A_DOUT({nc19860, nc19861, nc19862, nc19863, nc19864, nc19865, 
        nc19866, nc19867, nc19868, nc19869, nc19870, nc19871, nc19872, 
        nc19873, nc19874, \A_DOUT_TEMPR18[39] , \A_DOUT_TEMPR18[38] , 
        \A_DOUT_TEMPR18[37] , \A_DOUT_TEMPR18[36] , 
        \A_DOUT_TEMPR18[35] }), .B_DOUT({nc19875, nc19876, nc19877, 
        nc19878, nc19879, nc19880, nc19881, nc19882, nc19883, nc19884, 
        nc19885, nc19886, nc19887, nc19888, nc19889, 
        \B_DOUT_TEMPR18[39] , \B_DOUT_TEMPR18[38] , 
        \B_DOUT_TEMPR18[37] , \B_DOUT_TEMPR18[36] , 
        \B_DOUT_TEMPR18[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2622 (.A(\A_DOUT_TEMPR20[5] ), .B(\A_DOUT_TEMPR21[5] ), .C(
        \A_DOUT_TEMPR22[5] ), .D(\A_DOUT_TEMPR23[5] ), .Y(OR4_2622_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%93%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R93C3 (
        .A_DOUT({nc19890, nc19891, nc19892, nc19893, nc19894, nc19895, 
        nc19896, nc19897, nc19898, nc19899, nc19900, nc19901, nc19902, 
        nc19903, nc19904, \A_DOUT_TEMPR93[19] , \A_DOUT_TEMPR93[18] , 
        \A_DOUT_TEMPR93[17] , \A_DOUT_TEMPR93[16] , 
        \A_DOUT_TEMPR93[15] }), .B_DOUT({nc19905, nc19906, nc19907, 
        nc19908, nc19909, nc19910, nc19911, nc19912, nc19913, nc19914, 
        nc19915, nc19916, nc19917, nc19918, nc19919, 
        \B_DOUT_TEMPR93[19] , \B_DOUT_TEMPR93[18] , 
        \B_DOUT_TEMPR93[17] , \B_DOUT_TEMPR93[16] , 
        \B_DOUT_TEMPR93[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[93][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_857 (.A(OR4_2094_Y), .B(OR4_2467_Y), .C(OR4_68_Y), .D(
        OR4_2279_Y), .Y(OR4_857_Y));
    OR4 OR4_2978 (.A(\B_DOUT_TEMPR0[8] ), .B(\B_DOUT_TEMPR1[8] ), .C(
        \B_DOUT_TEMPR2[8] ), .D(\B_DOUT_TEMPR3[8] ), .Y(OR4_2978_Y));
    OR4 OR4_2285 (.A(\B_DOUT_TEMPR60[1] ), .B(\B_DOUT_TEMPR61[1] ), .C(
        \B_DOUT_TEMPR62[1] ), .D(\B_DOUT_TEMPR63[1] ), .Y(OR4_2285_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%87%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R87C0 (
        .A_DOUT({nc19920, nc19921, nc19922, nc19923, nc19924, nc19925, 
        nc19926, nc19927, nc19928, nc19929, nc19930, nc19931, nc19932, 
        nc19933, nc19934, \A_DOUT_TEMPR87[4] , \A_DOUT_TEMPR87[3] , 
        \A_DOUT_TEMPR87[2] , \A_DOUT_TEMPR87[1] , \A_DOUT_TEMPR87[0] })
        , .B_DOUT({nc19935, nc19936, nc19937, nc19938, nc19939, 
        nc19940, nc19941, nc19942, nc19943, nc19944, nc19945, nc19946, 
        nc19947, nc19948, nc19949, \B_DOUT_TEMPR87[4] , 
        \B_DOUT_TEMPR87[3] , \B_DOUT_TEMPR87[2] , \B_DOUT_TEMPR87[1] , 
        \B_DOUT_TEMPR87[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[87][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%95%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R95C3 (
        .A_DOUT({nc19950, nc19951, nc19952, nc19953, nc19954, nc19955, 
        nc19956, nc19957, nc19958, nc19959, nc19960, nc19961, nc19962, 
        nc19963, nc19964, \A_DOUT_TEMPR95[19] , \A_DOUT_TEMPR95[18] , 
        \A_DOUT_TEMPR95[17] , \A_DOUT_TEMPR95[16] , 
        \A_DOUT_TEMPR95[15] }), .B_DOUT({nc19965, nc19966, nc19967, 
        nc19968, nc19969, nc19970, nc19971, nc19972, nc19973, nc19974, 
        nc19975, nc19976, nc19977, nc19978, nc19979, 
        \B_DOUT_TEMPR95[19] , \B_DOUT_TEMPR95[18] , 
        \B_DOUT_TEMPR95[17] , \B_DOUT_TEMPR95[16] , 
        \B_DOUT_TEMPR95[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[95][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2907 (.A(\B_DOUT_TEMPR24[15] ), .B(\B_DOUT_TEMPR25[15] ), 
        .C(\B_DOUT_TEMPR26[15] ), .D(\B_DOUT_TEMPR27[15] ), .Y(
        OR4_2907_Y));
    OR4 OR4_1142 (.A(OR4_470_Y), .B(OR4_1413_Y), .C(OR4_2096_Y), .D(
        OR4_2392_Y), .Y(OR4_1142_Y));
    OR4 OR4_1425 (.A(OR4_622_Y), .B(OR4_2608_Y), .C(OR4_1238_Y), .D(
        OR4_2181_Y), .Y(OR4_1425_Y));
    OR4 OR4_2922 (.A(\A_DOUT_TEMPR79[39] ), .B(\A_DOUT_TEMPR80[39] ), 
        .C(\A_DOUT_TEMPR81[39] ), .D(\A_DOUT_TEMPR82[39] ), .Y(
        OR4_2922_Y));
    OR4 \OR4_B_DOUT[29]  (.A(OR4_387_Y), .B(OR4_1716_Y), .C(OR4_374_Y), 
        .D(OR4_2214_Y), .Y(B_DOUT[29]));
    OR4 OR4_1219 (.A(OR4_2434_Y), .B(OR4_308_Y), .C(OR4_3022_Y), .D(
        OR4_1457_Y), .Y(OR4_1219_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%33%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R33C2 (
        .A_DOUT({nc19980, nc19981, nc19982, nc19983, nc19984, nc19985, 
        nc19986, nc19987, nc19988, nc19989, nc19990, nc19991, nc19992, 
        nc19993, nc19994, \A_DOUT_TEMPR33[14] , \A_DOUT_TEMPR33[13] , 
        \A_DOUT_TEMPR33[12] , \A_DOUT_TEMPR33[11] , 
        \A_DOUT_TEMPR33[10] }), .B_DOUT({nc19995, nc19996, nc19997, 
        nc19998, nc19999, nc20000, nc20001, nc20002, nc20003, nc20004, 
        nc20005, nc20006, nc20007, nc20008, nc20009, 
        \B_DOUT_TEMPR33[14] , \B_DOUT_TEMPR33[13] , 
        \B_DOUT_TEMPR33[12] , \B_DOUT_TEMPR33[11] , 
        \B_DOUT_TEMPR33[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[33][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_76 (.A(\B_DOUT_TEMPR115[17] ), .B(\B_DOUT_TEMPR116[17] ), 
        .C(\B_DOUT_TEMPR117[17] ), .D(\B_DOUT_TEMPR118[17] ), .Y(
        OR4_76_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%27%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R27C4 (
        .A_DOUT({nc20010, nc20011, nc20012, nc20013, nc20014, nc20015, 
        nc20016, nc20017, nc20018, nc20019, nc20020, nc20021, nc20022, 
        nc20023, nc20024, \A_DOUT_TEMPR27[24] , \A_DOUT_TEMPR27[23] , 
        \A_DOUT_TEMPR27[22] , \A_DOUT_TEMPR27[21] , 
        \A_DOUT_TEMPR27[20] }), .B_DOUT({nc20025, nc20026, nc20027, 
        nc20028, nc20029, nc20030, nc20031, nc20032, nc20033, nc20034, 
        nc20035, nc20036, nc20037, nc20038, nc20039, 
        \B_DOUT_TEMPR27[24] , \B_DOUT_TEMPR27[23] , 
        \B_DOUT_TEMPR27[22] , \B_DOUT_TEMPR27[21] , 
        \B_DOUT_TEMPR27[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[27][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1470 (.A(OR4_869_Y), .B(OR4_669_Y), .C(OR2_18_Y), .D(
        \B_DOUT_TEMPR74[31] ), .Y(OR4_1470_Y));
    OR4 OR4_1958 (.A(\A_DOUT_TEMPR91[2] ), .B(\A_DOUT_TEMPR92[2] ), .C(
        \A_DOUT_TEMPR93[2] ), .D(\A_DOUT_TEMPR94[2] ), .Y(OR4_1958_Y));
    OR4 OR4_2364 (.A(\B_DOUT_TEMPR115[7] ), .B(\B_DOUT_TEMPR116[7] ), 
        .C(\B_DOUT_TEMPR117[7] ), .D(\B_DOUT_TEMPR118[7] ), .Y(
        OR4_2364_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%103%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R103C0 (
        .A_DOUT({nc20040, nc20041, nc20042, nc20043, nc20044, nc20045, 
        nc20046, nc20047, nc20048, nc20049, nc20050, nc20051, nc20052, 
        nc20053, nc20054, \A_DOUT_TEMPR103[4] , \A_DOUT_TEMPR103[3] , 
        \A_DOUT_TEMPR103[2] , \A_DOUT_TEMPR103[1] , 
        \A_DOUT_TEMPR103[0] }), .B_DOUT({nc20055, nc20056, nc20057, 
        nc20058, nc20059, nc20060, nc20061, nc20062, nc20063, nc20064, 
        nc20065, nc20066, nc20067, nc20068, nc20069, 
        \B_DOUT_TEMPR103[4] , \B_DOUT_TEMPR103[3] , 
        \B_DOUT_TEMPR103[2] , \B_DOUT_TEMPR103[1] , 
        \B_DOUT_TEMPR103[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[103][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1668 (.A(\B_DOUT_TEMPR36[28] ), .B(\B_DOUT_TEMPR37[28] ), 
        .C(\B_DOUT_TEMPR38[28] ), .D(\B_DOUT_TEMPR39[28] ), .Y(
        OR4_1668_Y));
    OR4 OR4_624 (.A(OR4_2862_Y), .B(OR4_2657_Y), .C(OR4_2606_Y), .D(
        OR4_512_Y), .Y(OR4_624_Y));
    OR4 OR4_2234 (.A(\A_DOUT_TEMPR99[35] ), .B(\A_DOUT_TEMPR100[35] ), 
        .C(\A_DOUT_TEMPR101[35] ), .D(\A_DOUT_TEMPR102[35] ), .Y(
        OR4_2234_Y));
    OR4 OR4_1489 (.A(\A_DOUT_TEMPR8[32] ), .B(\A_DOUT_TEMPR9[32] ), .C(
        \A_DOUT_TEMPR10[32] ), .D(\A_DOUT_TEMPR11[32] ), .Y(OR4_1489_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%1%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R1C0 (
        .A_DOUT({nc20070, nc20071, nc20072, nc20073, nc20074, nc20075, 
        nc20076, nc20077, nc20078, nc20079, nc20080, nc20081, nc20082, 
        nc20083, nc20084, \A_DOUT_TEMPR1[4] , \A_DOUT_TEMPR1[3] , 
        \A_DOUT_TEMPR1[2] , \A_DOUT_TEMPR1[1] , \A_DOUT_TEMPR1[0] }), 
        .B_DOUT({nc20085, nc20086, nc20087, nc20088, nc20089, nc20090, 
        nc20091, nc20092, nc20093, nc20094, nc20095, nc20096, nc20097, 
        nc20098, nc20099, \B_DOUT_TEMPR1[4] , \B_DOUT_TEMPR1[3] , 
        \B_DOUT_TEMPR1[2] , \B_DOUT_TEMPR1[1] , \B_DOUT_TEMPR1[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[1][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[0] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[0] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%75%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R75C7 (
        .A_DOUT({nc20100, nc20101, nc20102, nc20103, nc20104, nc20105, 
        nc20106, nc20107, nc20108, nc20109, nc20110, nc20111, nc20112, 
        nc20113, nc20114, \A_DOUT_TEMPR75[39] , \A_DOUT_TEMPR75[38] , 
        \A_DOUT_TEMPR75[37] , \A_DOUT_TEMPR75[36] , 
        \A_DOUT_TEMPR75[35] }), .B_DOUT({nc20115, nc20116, nc20117, 
        nc20118, nc20119, nc20120, nc20121, nc20122, nc20123, nc20124, 
        nc20125, nc20126, nc20127, nc20128, nc20129, 
        \B_DOUT_TEMPR75[39] , \B_DOUT_TEMPR75[38] , 
        \B_DOUT_TEMPR75[37] , \B_DOUT_TEMPR75[36] , 
        \B_DOUT_TEMPR75[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[75][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1726 (.A(\B_DOUT_TEMPR0[37] ), .B(\B_DOUT_TEMPR1[37] ), .C(
        \B_DOUT_TEMPR2[37] ), .D(\B_DOUT_TEMPR3[37] ), .Y(OR4_1726_Y));
    OR4 OR4_2800 (.A(\B_DOUT_TEMPR107[36] ), .B(\B_DOUT_TEMPR108[36] ), 
        .C(\B_DOUT_TEMPR109[36] ), .D(\B_DOUT_TEMPR110[36] ), .Y(
        OR4_2800_Y));
    OR2 OR2_53 (.A(\B_DOUT_TEMPR72[36] ), .B(\B_DOUT_TEMPR73[36] ), .Y(
        OR2_53_Y));
    OR4 OR4_1234 (.A(\B_DOUT_TEMPR4[25] ), .B(\B_DOUT_TEMPR5[25] ), .C(
        \B_DOUT_TEMPR6[25] ), .D(\B_DOUT_TEMPR7[25] ), .Y(OR4_1234_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%90%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R90C1 (
        .A_DOUT({nc20130, nc20131, nc20132, nc20133, nc20134, nc20135, 
        nc20136, nc20137, nc20138, nc20139, nc20140, nc20141, nc20142, 
        nc20143, nc20144, \A_DOUT_TEMPR90[9] , \A_DOUT_TEMPR90[8] , 
        \A_DOUT_TEMPR90[7] , \A_DOUT_TEMPR90[6] , \A_DOUT_TEMPR90[5] })
        , .B_DOUT({nc20145, nc20146, nc20147, nc20148, nc20149, 
        nc20150, nc20151, nc20152, nc20153, nc20154, nc20155, nc20156, 
        nc20157, nc20158, nc20159, \B_DOUT_TEMPR90[9] , 
        \B_DOUT_TEMPR90[8] , \B_DOUT_TEMPR90[7] , \B_DOUT_TEMPR90[6] , 
        \B_DOUT_TEMPR90[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[90][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2177 (.A(\A_DOUT_TEMPR4[23] ), .B(\A_DOUT_TEMPR5[23] ), .C(
        \A_DOUT_TEMPR6[23] ), .D(\A_DOUT_TEMPR7[23] ), .Y(OR4_2177_Y));
    OR4 OR4_1275 (.A(\A_DOUT_TEMPR79[26] ), .B(\A_DOUT_TEMPR80[26] ), 
        .C(\A_DOUT_TEMPR81[26] ), .D(\A_DOUT_TEMPR82[26] ), .Y(
        OR4_1275_Y));
    OR4 OR4_2674 (.A(\A_DOUT_TEMPR68[20] ), .B(\A_DOUT_TEMPR69[20] ), 
        .C(\A_DOUT_TEMPR70[20] ), .D(\A_DOUT_TEMPR71[20] ), .Y(
        OR4_2674_Y));
    OR4 OR4_2259 (.A(OR4_191_Y), .B(OR4_1398_Y), .C(OR2_60_Y), .D(
        \B_DOUT_TEMPR74[12] ), .Y(OR4_2259_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%23%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R23C6 (
        .A_DOUT({nc20160, nc20161, nc20162, nc20163, nc20164, nc20165, 
        nc20166, nc20167, nc20168, nc20169, nc20170, nc20171, nc20172, 
        nc20173, nc20174, \A_DOUT_TEMPR23[34] , \A_DOUT_TEMPR23[33] , 
        \A_DOUT_TEMPR23[32] , \A_DOUT_TEMPR23[31] , 
        \A_DOUT_TEMPR23[30] }), .B_DOUT({nc20175, nc20176, nc20177, 
        nc20178, nc20179, nc20180, nc20181, nc20182, nc20183, nc20184, 
        nc20185, nc20186, nc20187, nc20188, nc20189, 
        \B_DOUT_TEMPR23[34] , \B_DOUT_TEMPR23[33] , 
        \B_DOUT_TEMPR23[32] , \B_DOUT_TEMPR23[31] , 
        \B_DOUT_TEMPR23[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2696 (.A(\A_DOUT_TEMPR68[30] ), .B(\A_DOUT_TEMPR69[30] ), 
        .C(\A_DOUT_TEMPR70[30] ), .D(\A_DOUT_TEMPR71[30] ), .Y(
        OR4_2696_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%39%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R39C4 (
        .A_DOUT({nc20190, nc20191, nc20192, nc20193, nc20194, nc20195, 
        nc20196, nc20197, nc20198, nc20199, nc20200, nc20201, nc20202, 
        nc20203, nc20204, \A_DOUT_TEMPR39[24] , \A_DOUT_TEMPR39[23] , 
        \A_DOUT_TEMPR39[22] , \A_DOUT_TEMPR39[21] , 
        \A_DOUT_TEMPR39[20] }), .B_DOUT({nc20205, nc20206, nc20207, 
        nc20208, nc20209, nc20210, nc20211, nc20212, nc20213, nc20214, 
        nc20215, nc20216, nc20217, nc20218, nc20219, 
        \B_DOUT_TEMPR39[24] , \B_DOUT_TEMPR39[23] , 
        \B_DOUT_TEMPR39[22] , \B_DOUT_TEMPR39[21] , 
        \B_DOUT_TEMPR39[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[39][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_879 (.A(\A_DOUT_TEMPR95[28] ), .B(\A_DOUT_TEMPR96[28] ), 
        .C(\A_DOUT_TEMPR97[28] ), .D(\A_DOUT_TEMPR98[28] ), .Y(
        OR4_879_Y));
    OR4 OR4_2804 (.A(OR4_1421_Y), .B(OR4_1695_Y), .C(OR4_1202_Y), .D(
        OR4_2253_Y), .Y(OR4_2804_Y));
    OR4 OR4_2033 (.A(\A_DOUT_TEMPR115[16] ), .B(\A_DOUT_TEMPR116[16] ), 
        .C(\A_DOUT_TEMPR117[16] ), .D(\A_DOUT_TEMPR118[16] ), .Y(
        OR4_2033_Y));
    OR4 OR4_2190 (.A(\A_DOUT_TEMPR87[16] ), .B(\A_DOUT_TEMPR88[16] ), 
        .C(\A_DOUT_TEMPR89[16] ), .D(\A_DOUT_TEMPR90[16] ), .Y(
        OR4_2190_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%11%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R11C1 (
        .A_DOUT({nc20220, nc20221, nc20222, nc20223, nc20224, nc20225, 
        nc20226, nc20227, nc20228, nc20229, nc20230, nc20231, nc20232, 
        nc20233, nc20234, \A_DOUT_TEMPR11[9] , \A_DOUT_TEMPR11[8] , 
        \A_DOUT_TEMPR11[7] , \A_DOUT_TEMPR11[6] , \A_DOUT_TEMPR11[5] })
        , .B_DOUT({nc20235, nc20236, nc20237, nc20238, nc20239, 
        nc20240, nc20241, nc20242, nc20243, nc20244, nc20245, nc20246, 
        nc20247, nc20248, nc20249, \B_DOUT_TEMPR11[9] , 
        \B_DOUT_TEMPR11[8] , \B_DOUT_TEMPR11[7] , \B_DOUT_TEMPR11[6] , 
        \B_DOUT_TEMPR11[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_3013 (.A(OR4_1396_Y), .B(OR4_1139_Y), .C(OR4_1170_Y), .D(
        OR4_721_Y), .Y(OR4_3013_Y));
    OR4 OR4_2631 (.A(\A_DOUT_TEMPR44[11] ), .B(\A_DOUT_TEMPR45[11] ), 
        .C(\A_DOUT_TEMPR46[11] ), .D(\A_DOUT_TEMPR47[11] ), .Y(
        OR4_2631_Y));
    OR4 OR4_1033 (.A(\B_DOUT_TEMPR48[4] ), .B(\B_DOUT_TEMPR49[4] ), .C(
        \B_DOUT_TEMPR50[4] ), .D(\B_DOUT_TEMPR51[4] ), .Y(OR4_1033_Y));
    OR4 OR4_271 (.A(\A_DOUT_TEMPR75[17] ), .B(\A_DOUT_TEMPR76[17] ), 
        .C(\A_DOUT_TEMPR77[17] ), .D(\A_DOUT_TEMPR78[17] ), .Y(
        OR4_271_Y));
    OR4 OR4_1380 (.A(OR4_715_Y), .B(OR4_1713_Y), .C(OR4_1216_Y), .D(
        OR4_1559_Y), .Y(OR4_1380_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%112%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R112C1 (
        .A_DOUT({nc20250, nc20251, nc20252, nc20253, nc20254, nc20255, 
        nc20256, nc20257, nc20258, nc20259, nc20260, nc20261, nc20262, 
        nc20263, nc20264, \A_DOUT_TEMPR112[9] , \A_DOUT_TEMPR112[8] , 
        \A_DOUT_TEMPR112[7] , \A_DOUT_TEMPR112[6] , 
        \A_DOUT_TEMPR112[5] }), .B_DOUT({nc20265, nc20266, nc20267, 
        nc20268, nc20269, nc20270, nc20271, nc20272, nc20273, nc20274, 
        nc20275, nc20276, nc20277, nc20278, nc20279, 
        \B_DOUT_TEMPR112[9] , \B_DOUT_TEMPR112[8] , 
        \B_DOUT_TEMPR112[7] , \B_DOUT_TEMPR112[6] , 
        \B_DOUT_TEMPR112[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[112][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_871 (.A(\B_DOUT_TEMPR52[10] ), .B(\B_DOUT_TEMPR53[10] ), 
        .C(\B_DOUT_TEMPR54[10] ), .D(\B_DOUT_TEMPR55[10] ), .Y(
        OR4_871_Y));
    OR4 OR4_1592 (.A(\A_DOUT_TEMPR107[15] ), .B(\A_DOUT_TEMPR108[15] ), 
        .C(\A_DOUT_TEMPR109[15] ), .D(\A_DOUT_TEMPR110[15] ), .Y(
        OR4_1592_Y));
    OR4 OR4_1487 (.A(\B_DOUT_TEMPR44[28] ), .B(\B_DOUT_TEMPR45[28] ), 
        .C(\B_DOUT_TEMPR46[28] ), .D(\B_DOUT_TEMPR47[28] ), .Y(
        OR4_1487_Y));
    OR4 OR4_632 (.A(\A_DOUT_TEMPR52[19] ), .B(\A_DOUT_TEMPR53[19] ), 
        .C(\A_DOUT_TEMPR54[19] ), .D(\A_DOUT_TEMPR55[19] ), .Y(
        OR4_632_Y));
    OR4 OR4_2733 (.A(\A_DOUT_TEMPR36[5] ), .B(\A_DOUT_TEMPR37[5] ), .C(
        \A_DOUT_TEMPR38[5] ), .D(\A_DOUT_TEMPR39[5] ), .Y(OR4_2733_Y));
    OR4 OR4_1157 (.A(\B_DOUT_TEMPR12[10] ), .B(\B_DOUT_TEMPR13[10] ), 
        .C(\B_DOUT_TEMPR14[10] ), .D(\B_DOUT_TEMPR15[10] ), .Y(
        OR4_1157_Y));
    OR4 OR4_1631 (.A(\A_DOUT_TEMPR4[25] ), .B(\A_DOUT_TEMPR5[25] ), .C(
        \A_DOUT_TEMPR6[25] ), .D(\A_DOUT_TEMPR7[25] ), .Y(OR4_1631_Y));
    OR4 OR4_1654 (.A(\A_DOUT_TEMPR24[20] ), .B(\A_DOUT_TEMPR25[20] ), 
        .C(\A_DOUT_TEMPR26[20] ), .D(\A_DOUT_TEMPR27[20] ), .Y(
        OR4_1654_Y));
    OR2 OR2_41 (.A(\A_DOUT_TEMPR72[15] ), .B(\A_DOUT_TEMPR73[15] ), .Y(
        OR2_41_Y));
    OR4 OR4_67 (.A(\B_DOUT_TEMPR12[26] ), .B(\B_DOUT_TEMPR13[26] ), .C(
        \B_DOUT_TEMPR14[26] ), .D(\B_DOUT_TEMPR15[26] ), .Y(OR4_67_Y));
    OR4 OR4_2135 (.A(\B_DOUT_TEMPR4[15] ), .B(\B_DOUT_TEMPR5[15] ), .C(
        \B_DOUT_TEMPR6[15] ), .D(\B_DOUT_TEMPR7[15] ), .Y(OR4_2135_Y));
    OR4 OR4_1733 (.A(\A_DOUT_TEMPR36[15] ), .B(\A_DOUT_TEMPR37[15] ), 
        .C(\A_DOUT_TEMPR38[15] ), .D(\A_DOUT_TEMPR39[15] ), .Y(
        OR4_1733_Y));
    OR4 OR4_2429 (.A(\B_DOUT_TEMPR68[32] ), .B(\B_DOUT_TEMPR69[32] ), 
        .C(\B_DOUT_TEMPR70[32] ), .D(\B_DOUT_TEMPR71[32] ), .Y(
        OR4_2429_Y));
    OR4 OR4_2686 (.A(\B_DOUT_TEMPR8[35] ), .B(\B_DOUT_TEMPR9[35] ), .C(
        \B_DOUT_TEMPR10[35] ), .D(\B_DOUT_TEMPR11[35] ), .Y(OR4_2686_Y)
        );
    OR4 OR4_1135 (.A(\A_DOUT_TEMPR111[39] ), .B(\A_DOUT_TEMPR112[39] ), 
        .C(\A_DOUT_TEMPR113[39] ), .D(\A_DOUT_TEMPR114[39] ), .Y(
        OR4_1135_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%105%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R105C7 (
        .A_DOUT({nc20280, nc20281, nc20282, nc20283, nc20284, nc20285, 
        nc20286, nc20287, nc20288, nc20289, nc20290, nc20291, nc20292, 
        nc20293, nc20294, \A_DOUT_TEMPR105[39] , \A_DOUT_TEMPR105[38] , 
        \A_DOUT_TEMPR105[37] , \A_DOUT_TEMPR105[36] , 
        \A_DOUT_TEMPR105[35] }), .B_DOUT({nc20295, nc20296, nc20297, 
        nc20298, nc20299, nc20300, nc20301, nc20302, nc20303, nc20304, 
        nc20305, nc20306, nc20307, nc20308, nc20309, 
        \B_DOUT_TEMPR105[39] , \B_DOUT_TEMPR105[38] , 
        \B_DOUT_TEMPR105[37] , \B_DOUT_TEMPR105[36] , 
        \B_DOUT_TEMPR105[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[105][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_451 (.A(\A_DOUT_TEMPR87[9] ), .B(\A_DOUT_TEMPR88[9] ), .C(
        \A_DOUT_TEMPR89[9] ), .D(\A_DOUT_TEMPR90[9] ), .Y(OR4_451_Y));
    OR4 OR4_2180 (.A(\B_DOUT_TEMPR95[17] ), .B(\B_DOUT_TEMPR96[17] ), 
        .C(\B_DOUT_TEMPR97[17] ), .D(\B_DOUT_TEMPR98[17] ), .Y(
        OR4_2180_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%106%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R106C7 (
        .A_DOUT({nc20310, nc20311, nc20312, nc20313, nc20314, nc20315, 
        nc20316, nc20317, nc20318, nc20319, nc20320, nc20321, nc20322, 
        nc20323, nc20324, \A_DOUT_TEMPR106[39] , \A_DOUT_TEMPR106[38] , 
        \A_DOUT_TEMPR106[37] , \A_DOUT_TEMPR106[36] , 
        \A_DOUT_TEMPR106[35] }), .B_DOUT({nc20325, nc20326, nc20327, 
        nc20328, nc20329, nc20330, nc20331, nc20332, nc20333, nc20334, 
        nc20335, nc20336, nc20337, nc20338, nc20339, 
        \B_DOUT_TEMPR106[39] , \B_DOUT_TEMPR106[38] , 
        \B_DOUT_TEMPR106[37] , \B_DOUT_TEMPR106[36] , 
        \B_DOUT_TEMPR106[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[106][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%113%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R113C1 (
        .A_DOUT({nc20340, nc20341, nc20342, nc20343, nc20344, nc20345, 
        nc20346, nc20347, nc20348, nc20349, nc20350, nc20351, nc20352, 
        nc20353, nc20354, \A_DOUT_TEMPR113[9] , \A_DOUT_TEMPR113[8] , 
        \A_DOUT_TEMPR113[7] , \A_DOUT_TEMPR113[6] , 
        \A_DOUT_TEMPR113[5] }), .B_DOUT({nc20355, nc20356, nc20357, 
        nc20358, nc20359, nc20360, nc20361, nc20362, nc20363, nc20364, 
        nc20365, nc20366, nc20367, nc20368, nc20369, 
        \B_DOUT_TEMPR113[9] , \B_DOUT_TEMPR113[8] , 
        \B_DOUT_TEMPR113[7] , \B_DOUT_TEMPR113[6] , 
        \B_DOUT_TEMPR113[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[113][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2031 (.A(OR4_1597_Y), .B(OR4_2407_Y), .C(OR2_35_Y), .D(
        \B_DOUT_TEMPR74[22] ), .Y(OR4_2031_Y));
    OR4 OR4_644 (.A(\A_DOUT_TEMPR52[16] ), .B(\A_DOUT_TEMPR53[16] ), 
        .C(\A_DOUT_TEMPR54[16] ), .D(\A_DOUT_TEMPR55[16] ), .Y(
        OR4_644_Y));
    OR4 OR4_3011 (.A(\A_DOUT_TEMPR60[34] ), .B(\A_DOUT_TEMPR61[34] ), 
        .C(\A_DOUT_TEMPR62[34] ), .D(\A_DOUT_TEMPR63[34] ), .Y(
        OR4_3011_Y));
    OR4 OR4_897 (.A(\B_DOUT_TEMPR95[36] ), .B(\B_DOUT_TEMPR96[36] ), 
        .C(\B_DOUT_TEMPR97[36] ), .D(\B_DOUT_TEMPR98[36] ), .Y(
        OR4_897_Y));
    OR4 OR4_809 (.A(\B_DOUT_TEMPR87[22] ), .B(\B_DOUT_TEMPR88[22] ), 
        .C(\B_DOUT_TEMPR89[22] ), .D(\B_DOUT_TEMPR90[22] ), .Y(
        OR4_809_Y));
    OR4 OR4_2460 (.A(OR4_2854_Y), .B(OR4_161_Y), .C(OR4_949_Y), .D(
        OR4_1723_Y), .Y(OR4_2460_Y));
    OR4 OR4_1031 (.A(\A_DOUT_TEMPR0[10] ), .B(\A_DOUT_TEMPR1[10] ), .C(
        \A_DOUT_TEMPR2[10] ), .D(\A_DOUT_TEMPR3[10] ), .Y(OR4_1031_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%44%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R44C0 (
        .A_DOUT({nc20370, nc20371, nc20372, nc20373, nc20374, nc20375, 
        nc20376, nc20377, nc20378, nc20379, nc20380, nc20381, nc20382, 
        nc20383, nc20384, \A_DOUT_TEMPR44[4] , \A_DOUT_TEMPR44[3] , 
        \A_DOUT_TEMPR44[2] , \A_DOUT_TEMPR44[1] , \A_DOUT_TEMPR44[0] })
        , .B_DOUT({nc20385, nc20386, nc20387, nc20388, nc20389, 
        nc20390, nc20391, nc20392, nc20393, nc20394, nc20395, nc20396, 
        nc20397, nc20398, nc20399, \B_DOUT_TEMPR44[4] , 
        \B_DOUT_TEMPR44[3] , \B_DOUT_TEMPR44[2] , \B_DOUT_TEMPR44[1] , 
        \B_DOUT_TEMPR44[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[44][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1249 (.A(\A_DOUT_TEMPR20[4] ), .B(\A_DOUT_TEMPR21[4] ), .C(
        \A_DOUT_TEMPR22[4] ), .D(\A_DOUT_TEMPR23[4] ), .Y(OR4_1249_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%24%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R24C4 (
        .A_DOUT({nc20400, nc20401, nc20402, nc20403, nc20404, nc20405, 
        nc20406, nc20407, nc20408, nc20409, nc20410, nc20411, nc20412, 
        nc20413, nc20414, \A_DOUT_TEMPR24[24] , \A_DOUT_TEMPR24[23] , 
        \A_DOUT_TEMPR24[22] , \A_DOUT_TEMPR24[21] , 
        \A_DOUT_TEMPR24[20] }), .B_DOUT({nc20415, nc20416, nc20417, 
        nc20418, nc20419, nc20420, nc20421, nc20422, nc20423, nc20424, 
        nc20425, nc20426, nc20427, nc20428, nc20429, 
        \B_DOUT_TEMPR24[24] , \B_DOUT_TEMPR24[23] , 
        \B_DOUT_TEMPR24[22] , \B_DOUT_TEMPR24[21] , 
        \B_DOUT_TEMPR24[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2320 (.A(\A_DOUT_TEMPR111[12] ), .B(\A_DOUT_TEMPR112[12] ), 
        .C(\A_DOUT_TEMPR113[12] ), .D(\A_DOUT_TEMPR114[12] ), .Y(
        OR4_2320_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%89%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R89C6 (
        .A_DOUT({nc20430, nc20431, nc20432, nc20433, nc20434, nc20435, 
        nc20436, nc20437, nc20438, nc20439, nc20440, nc20441, nc20442, 
        nc20443, nc20444, \A_DOUT_TEMPR89[34] , \A_DOUT_TEMPR89[33] , 
        \A_DOUT_TEMPR89[32] , \A_DOUT_TEMPR89[31] , 
        \A_DOUT_TEMPR89[30] }), .B_DOUT({nc20445, nc20446, nc20447, 
        nc20448, nc20449, nc20450, nc20451, nc20452, nc20453, nc20454, 
        nc20455, nc20456, nc20457, nc20458, nc20459, 
        \B_DOUT_TEMPR89[34] , \B_DOUT_TEMPR89[33] , 
        \B_DOUT_TEMPR89[32] , \B_DOUT_TEMPR89[31] , 
        \B_DOUT_TEMPR89[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[89][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2427 (.A(OR4_594_Y), .B(OR4_398_Y), .C(OR2_10_Y), .D(
        \B_DOUT_TEMPR74[39] ), .Y(OR4_2427_Y));
    OR4 OR4_466 (.A(\B_DOUT_TEMPR0[24] ), .B(\B_DOUT_TEMPR1[24] ), .C(
        \B_DOUT_TEMPR2[24] ), .D(\B_DOUT_TEMPR3[24] ), .Y(OR4_466_Y));
    OR4 OR4_201 (.A(\A_DOUT_TEMPR111[10] ), .B(\A_DOUT_TEMPR112[10] ), 
        .C(\A_DOUT_TEMPR113[10] ), .D(\A_DOUT_TEMPR114[10] ), .Y(
        OR4_201_Y));
    OR4 OR4_801 (.A(\A_DOUT_TEMPR87[30] ), .B(\A_DOUT_TEMPR88[30] ), 
        .C(\A_DOUT_TEMPR89[30] ), .D(\A_DOUT_TEMPR90[30] ), .Y(
        OR4_801_Y));
    OR4 OR4_627 (.A(\B_DOUT_TEMPR87[16] ), .B(\B_DOUT_TEMPR88[16] ), 
        .C(\B_DOUT_TEMPR89[16] ), .D(\B_DOUT_TEMPR90[16] ), .Y(
        OR4_627_Y));
    OR4 OR4_377 (.A(\B_DOUT_TEMPR12[12] ), .B(\B_DOUT_TEMPR13[12] ), 
        .C(\B_DOUT_TEMPR14[12] ), .D(\B_DOUT_TEMPR15[12] ), .Y(
        OR4_377_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%77%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R77C2 (
        .A_DOUT({nc20460, nc20461, nc20462, nc20463, nc20464, nc20465, 
        nc20466, nc20467, nc20468, nc20469, nc20470, nc20471, nc20472, 
        nc20473, nc20474, \A_DOUT_TEMPR77[14] , \A_DOUT_TEMPR77[13] , 
        \A_DOUT_TEMPR77[12] , \A_DOUT_TEMPR77[11] , 
        \A_DOUT_TEMPR77[10] }), .B_DOUT({nc20475, nc20476, nc20477, 
        nc20478, nc20479, nc20480, nc20481, nc20482, nc20483, nc20484, 
        nc20485, nc20486, nc20487, nc20488, nc20489, 
        \B_DOUT_TEMPR77[14] , \B_DOUT_TEMPR77[13] , 
        \B_DOUT_TEMPR77[12] , \B_DOUT_TEMPR77[11] , 
        \B_DOUT_TEMPR77[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[77][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_60 (.A(\A_DOUT_TEMPR28[0] ), .B(\A_DOUT_TEMPR29[0] ), .C(
        \A_DOUT_TEMPR30[0] ), .D(\A_DOUT_TEMPR31[0] ), .Y(OR4_60_Y));
    OR4 OR4_1676 (.A(\A_DOUT_TEMPR111[25] ), .B(\A_DOUT_TEMPR112[25] ), 
        .C(\A_DOUT_TEMPR113[25] ), .D(\A_DOUT_TEMPR114[25] ), .Y(
        OR4_1676_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%8%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R8C1 (
        .A_DOUT({nc20490, nc20491, nc20492, nc20493, nc20494, nc20495, 
        nc20496, nc20497, nc20498, nc20499, nc20500, nc20501, nc20502, 
        nc20503, nc20504, \A_DOUT_TEMPR8[9] , \A_DOUT_TEMPR8[8] , 
        \A_DOUT_TEMPR8[7] , \A_DOUT_TEMPR8[6] , \A_DOUT_TEMPR8[5] }), 
        .B_DOUT({nc20505, nc20506, nc20507, nc20508, nc20509, nc20510, 
        nc20511, nc20512, nc20513, nc20514, nc20515, nc20516, nc20517, 
        nc20518, nc20519, \B_DOUT_TEMPR8[9] , \B_DOUT_TEMPR8[8] , 
        \B_DOUT_TEMPR8[7] , \B_DOUT_TEMPR8[6] , \B_DOUT_TEMPR8[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[8][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[2] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1090 (.A(\B_DOUT_TEMPR4[35] ), .B(\B_DOUT_TEMPR5[35] ), .C(
        \B_DOUT_TEMPR6[35] ), .D(\B_DOUT_TEMPR7[35] ), .Y(OR4_1090_Y));
    OR4 OR4_878 (.A(\A_DOUT_TEMPR95[5] ), .B(\A_DOUT_TEMPR96[5] ), .C(
        \A_DOUT_TEMPR97[5] ), .D(\A_DOUT_TEMPR98[5] ), .Y(OR4_878_Y));
    OR4 OR4_1701 (.A(OR4_1206_Y), .B(OR4_1478_Y), .C(OR4_53_Y), .D(
        OR4_986_Y), .Y(OR4_1701_Y));
    OR4 OR4_2265 (.A(OR4_844_Y), .B(OR4_1978_Y), .C(OR4_2330_Y), .D(
        OR4_2666_Y), .Y(OR4_2265_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%46%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R46C7 (
        .A_DOUT({nc20520, nc20521, nc20522, nc20523, nc20524, nc20525, 
        nc20526, nc20527, nc20528, nc20529, nc20530, nc20531, nc20532, 
        nc20533, nc20534, \A_DOUT_TEMPR46[39] , \A_DOUT_TEMPR46[38] , 
        \A_DOUT_TEMPR46[37] , \A_DOUT_TEMPR46[36] , 
        \A_DOUT_TEMPR46[35] }), .B_DOUT({nc20535, nc20536, nc20537, 
        nc20538, nc20539, nc20540, nc20541, nc20542, nc20543, nc20544, 
        nc20545, nc20546, nc20547, nc20548, nc20549, 
        \B_DOUT_TEMPR46[39] , \B_DOUT_TEMPR46[38] , 
        \B_DOUT_TEMPR46[37] , \B_DOUT_TEMPR46[36] , 
        \B_DOUT_TEMPR46[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[46][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1170 (.A(OR4_1652_Y), .B(OR4_2396_Y), .C(OR4_860_Y), .D(
        OR4_2397_Y), .Y(OR4_1170_Y));
    OR4 OR4_671 (.A(\A_DOUT_TEMPR44[35] ), .B(\A_DOUT_TEMPR45[35] ), 
        .C(\A_DOUT_TEMPR46[35] ), .D(\A_DOUT_TEMPR47[35] ), .Y(
        OR4_671_Y));
    OR4 OR4_1527 (.A(\B_DOUT_TEMPR28[6] ), .B(\B_DOUT_TEMPR29[6] ), .C(
        \B_DOUT_TEMPR30[6] ), .D(\B_DOUT_TEMPR31[6] ), .Y(OR4_1527_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%63%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R63C2 (
        .A_DOUT({nc20550, nc20551, nc20552, nc20553, nc20554, nc20555, 
        nc20556, nc20557, nc20558, nc20559, nc20560, nc20561, nc20562, 
        nc20563, nc20564, \A_DOUT_TEMPR63[14] , \A_DOUT_TEMPR63[13] , 
        \A_DOUT_TEMPR63[12] , \A_DOUT_TEMPR63[11] , 
        \A_DOUT_TEMPR63[10] }), .B_DOUT({nc20565, nc20566, nc20567, 
        nc20568, nc20569, nc20570, nc20571, nc20572, nc20573, nc20574, 
        nc20575, nc20576, nc20577, nc20578, nc20579, 
        \B_DOUT_TEMPR63[14] , \B_DOUT_TEMPR63[13] , 
        \B_DOUT_TEMPR63[12] , \B_DOUT_TEMPR63[11] , 
        \B_DOUT_TEMPR63[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[63][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1869 (.A(\A_DOUT_TEMPR4[31] ), .B(\A_DOUT_TEMPR5[31] ), .C(
        \A_DOUT_TEMPR6[31] ), .D(\A_DOUT_TEMPR7[31] ), .Y(OR4_1869_Y));
    OR4 OR4_2993 (.A(\B_DOUT_TEMPR8[15] ), .B(\B_DOUT_TEMPR9[15] ), .C(
        \B_DOUT_TEMPR10[15] ), .D(\B_DOUT_TEMPR11[15] ), .Y(OR4_2993_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%47%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R47C6 (
        .A_DOUT({nc20580, nc20581, nc20582, nc20583, nc20584, nc20585, 
        nc20586, nc20587, nc20588, nc20589, nc20590, nc20591, nc20592, 
        nc20593, nc20594, \A_DOUT_TEMPR47[34] , \A_DOUT_TEMPR47[33] , 
        \A_DOUT_TEMPR47[32] , \A_DOUT_TEMPR47[31] , 
        \A_DOUT_TEMPR47[30] }), .B_DOUT({nc20595, nc20596, nc20597, 
        nc20598, nc20599, nc20600, nc20601, nc20602, nc20603, nc20604, 
        nc20605, nc20606, nc20607, nc20608, nc20609, 
        \B_DOUT_TEMPR47[34] , \B_DOUT_TEMPR47[33] , 
        \B_DOUT_TEMPR47[32] , \B_DOUT_TEMPR47[31] , 
        \B_DOUT_TEMPR47[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%53%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R53C3 (
        .A_DOUT({nc20610, nc20611, nc20612, nc20613, nc20614, nc20615, 
        nc20616, nc20617, nc20618, nc20619, nc20620, nc20621, nc20622, 
        nc20623, nc20624, \A_DOUT_TEMPR53[19] , \A_DOUT_TEMPR53[18] , 
        \A_DOUT_TEMPR53[17] , \A_DOUT_TEMPR53[16] , 
        \A_DOUT_TEMPR53[15] }), .B_DOUT({nc20625, nc20626, nc20627, 
        nc20628, nc20629, nc20630, nc20631, nc20632, nc20633, nc20634, 
        nc20635, nc20636, nc20637, nc20638, nc20639, 
        \B_DOUT_TEMPR53[19] , \B_DOUT_TEMPR53[18] , 
        \B_DOUT_TEMPR53[17] , \B_DOUT_TEMPR53[16] , 
        \B_DOUT_TEMPR53[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[53][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%90%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R90C7 (
        .A_DOUT({nc20640, nc20641, nc20642, nc20643, nc20644, nc20645, 
        nc20646, nc20647, nc20648, nc20649, nc20650, nc20651, nc20652, 
        nc20653, nc20654, \A_DOUT_TEMPR90[39] , \A_DOUT_TEMPR90[38] , 
        \A_DOUT_TEMPR90[37] , \A_DOUT_TEMPR90[36] , 
        \A_DOUT_TEMPR90[35] }), .B_DOUT({nc20655, nc20656, nc20657, 
        nc20658, nc20659, nc20660, nc20661, nc20662, nc20663, nc20664, 
        nc20665, nc20666, nc20667, nc20668, nc20669, 
        \B_DOUT_TEMPR90[39] , \B_DOUT_TEMPR90[38] , 
        \B_DOUT_TEMPR90[37] , \B_DOUT_TEMPR90[36] , 
        \B_DOUT_TEMPR90[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[90][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_47 (.A(\A_DOUT_TEMPR4[22] ), .B(\A_DOUT_TEMPR5[22] ), .C(
        \A_DOUT_TEMPR6[22] ), .D(\A_DOUT_TEMPR7[22] ), .Y(OR4_47_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%55%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R55C3 (
        .A_DOUT({nc20670, nc20671, nc20672, nc20673, nc20674, nc20675, 
        nc20676, nc20677, nc20678, nc20679, nc20680, nc20681, nc20682, 
        nc20683, nc20684, \A_DOUT_TEMPR55[19] , \A_DOUT_TEMPR55[18] , 
        \A_DOUT_TEMPR55[17] , \A_DOUT_TEMPR55[16] , 
        \A_DOUT_TEMPR55[15] }), .B_DOUT({nc20685, nc20686, nc20687, 
        nc20688, nc20689, nc20690, nc20691, nc20692, nc20693, nc20694, 
        nc20695, nc20696, nc20697, nc20698, nc20699, 
        \B_DOUT_TEMPR55[19] , \B_DOUT_TEMPR55[18] , 
        \B_DOUT_TEMPR55[17] , \B_DOUT_TEMPR55[16] , 
        \B_DOUT_TEMPR55[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[55][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2670 (.A(\A_DOUT_TEMPR52[2] ), .B(\A_DOUT_TEMPR53[2] ), .C(
        \A_DOUT_TEMPR54[2] ), .D(\A_DOUT_TEMPR55[2] ), .Y(OR4_2670_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENA[0]  (.A(A_WBYTE_EN[0]), .B(
        A_WEN), .Y(\WBYTEENA[0] ));
    OR4 OR4_1161 (.A(OR4_1612_Y), .B(OR4_644_Y), .C(OR4_858_Y), .D(
        OR4_659_Y), .Y(OR4_1161_Y));
    OR4 OR4_474 (.A(\B_DOUT_TEMPR56[22] ), .B(\B_DOUT_TEMPR57[22] ), 
        .C(\B_DOUT_TEMPR58[22] ), .D(\B_DOUT_TEMPR59[22] ), .Y(
        OR4_474_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%6%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R6C0 (
        .A_DOUT({nc20700, nc20701, nc20702, nc20703, nc20704, nc20705, 
        nc20706, nc20707, nc20708, nc20709, nc20710, nc20711, nc20712, 
        nc20713, nc20714, \A_DOUT_TEMPR6[4] , \A_DOUT_TEMPR6[3] , 
        \A_DOUT_TEMPR6[2] , \A_DOUT_TEMPR6[1] , \A_DOUT_TEMPR6[0] }), 
        .B_DOUT({nc20715, nc20716, nc20717, nc20718, nc20719, nc20720, 
        nc20721, nc20722, nc20723, nc20724, nc20725, nc20726, nc20727, 
        nc20728, nc20729, \B_DOUT_TEMPR6[4] , \B_DOUT_TEMPR6[3] , 
        \B_DOUT_TEMPR6[2] , \B_DOUT_TEMPR6[1] , \B_DOUT_TEMPR6[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[6][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[1] , A_ADDR[13], \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[1] , B_ADDR[13], \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2078 (.A(OR4_1906_Y), .B(OR4_2847_Y), .C(OR4_2463_Y), .D(
        OR4_958_Y), .Y(OR4_2078_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%42%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R42C4 (
        .A_DOUT({nc20730, nc20731, nc20732, nc20733, nc20734, nc20735, 
        nc20736, nc20737, nc20738, nc20739, nc20740, nc20741, nc20742, 
        nc20743, nc20744, \A_DOUT_TEMPR42[24] , \A_DOUT_TEMPR42[23] , 
        \A_DOUT_TEMPR42[22] , \A_DOUT_TEMPR42[21] , 
        \A_DOUT_TEMPR42[20] }), .B_DOUT({nc20745, nc20746, nc20747, 
        nc20748, nc20749, nc20750, nc20751, nc20752, nc20753, nc20754, 
        nc20755, nc20756, nc20757, nc20758, nc20759, 
        \B_DOUT_TEMPR42[24] , \B_DOUT_TEMPR42[23] , 
        \B_DOUT_TEMPR42[22] , \B_DOUT_TEMPR42[21] , 
        \B_DOUT_TEMPR42[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[42][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%87%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R87C1 (
        .A_DOUT({nc20760, nc20761, nc20762, nc20763, nc20764, nc20765, 
        nc20766, nc20767, nc20768, nc20769, nc20770, nc20771, nc20772, 
        nc20773, nc20774, \A_DOUT_TEMPR87[9] , \A_DOUT_TEMPR87[8] , 
        \A_DOUT_TEMPR87[7] , \A_DOUT_TEMPR87[6] , \A_DOUT_TEMPR87[5] })
        , .B_DOUT({nc20775, nc20776, nc20777, nc20778, nc20779, 
        nc20780, nc20781, nc20782, nc20783, nc20784, nc20785, nc20786, 
        nc20787, nc20788, nc20789, \B_DOUT_TEMPR87[9] , 
        \B_DOUT_TEMPR87[8] , \B_DOUT_TEMPR87[7] , \B_DOUT_TEMPR87[6] , 
        \B_DOUT_TEMPR87[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[87][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2305 (.A(\A_DOUT_TEMPR95[39] ), .B(\A_DOUT_TEMPR96[39] ), 
        .C(\A_DOUT_TEMPR97[39] ), .D(\A_DOUT_TEMPR98[39] ), .Y(
        OR4_2305_Y));
    OR4 OR4_227 (.A(\A_DOUT_TEMPR115[14] ), .B(\A_DOUT_TEMPR116[14] ), 
        .C(\A_DOUT_TEMPR117[14] ), .D(\A_DOUT_TEMPR118[14] ), .Y(
        OR4_227_Y));
    OR4 OR4_1065 (.A(\B_DOUT_TEMPR0[31] ), .B(\B_DOUT_TEMPR1[31] ), .C(
        \B_DOUT_TEMPR2[31] ), .D(\B_DOUT_TEMPR3[31] ), .Y(OR4_1065_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[11]  (.A(CFG3_20_Y), .B(
        CFG3_15_Y), .Y(\BLKY2[11] ));
    OR4 OR4_2391 (.A(\B_DOUT_TEMPR107[19] ), .B(\B_DOUT_TEMPR108[19] ), 
        .C(\B_DOUT_TEMPR109[19] ), .D(\B_DOUT_TEMPR110[19] ), .Y(
        OR4_2391_Y));
    OR4 OR4_210 (.A(\A_DOUT_TEMPR115[22] ), .B(\A_DOUT_TEMPR116[22] ), 
        .C(\A_DOUT_TEMPR117[22] ), .D(\A_DOUT_TEMPR118[22] ), .Y(
        OR4_210_Y));
    OR4 OR4_2983 (.A(\B_DOUT_TEMPR83[8] ), .B(\B_DOUT_TEMPR84[8] ), .C(
        \B_DOUT_TEMPR85[8] ), .D(\B_DOUT_TEMPR86[8] ), .Y(OR4_2983_Y));
    OR4 OR4_2891 (.A(\A_DOUT_TEMPR4[6] ), .B(\A_DOUT_TEMPR5[6] ), .C(
        \A_DOUT_TEMPR6[6] ), .D(\A_DOUT_TEMPR7[6] ), .Y(OR4_2891_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%69%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R69C4 (
        .A_DOUT({nc20790, nc20791, nc20792, nc20793, nc20794, nc20795, 
        nc20796, nc20797, nc20798, nc20799, nc20800, nc20801, nc20802, 
        nc20803, nc20804, \A_DOUT_TEMPR69[24] , \A_DOUT_TEMPR69[23] , 
        \A_DOUT_TEMPR69[22] , \A_DOUT_TEMPR69[21] , 
        \A_DOUT_TEMPR69[20] }), .B_DOUT({nc20805, nc20806, nc20807, 
        nc20808, nc20809, nc20810, nc20811, nc20812, nc20813, nc20814, 
        nc20815, nc20816, nc20817, nc20818, nc20819, 
        \B_DOUT_TEMPR69[24] , \B_DOUT_TEMPR69[23] , 
        \B_DOUT_TEMPR69[22] , \B_DOUT_TEMPR69[21] , 
        \B_DOUT_TEMPR69[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[69][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1650 (.A(\B_DOUT_TEMPR91[9] ), .B(\B_DOUT_TEMPR92[9] ), .C(
        \B_DOUT_TEMPR93[9] ), .D(\B_DOUT_TEMPR94[9] ), .Y(OR4_1650_Y));
    OR4 OR4_1911 (.A(\A_DOUT_TEMPR32[36] ), .B(\A_DOUT_TEMPR33[36] ), 
        .C(\A_DOUT_TEMPR34[36] ), .D(\A_DOUT_TEMPR35[36] ), .Y(
        OR4_1911_Y));
    OR4 OR4_307 (.A(\A_DOUT_TEMPR64[11] ), .B(\A_DOUT_TEMPR65[11] ), 
        .C(\A_DOUT_TEMPR66[11] ), .D(\A_DOUT_TEMPR67[11] ), .Y(
        OR4_307_Y));
    OR4 OR4_2142 (.A(\A_DOUT_TEMPR52[29] ), .B(\A_DOUT_TEMPR53[29] ), 
        .C(\A_DOUT_TEMPR54[29] ), .D(\A_DOUT_TEMPR55[29] ), .Y(
        OR4_2142_Y));
    OR4 OR4_610 (.A(\B_DOUT_TEMPR95[38] ), .B(\B_DOUT_TEMPR96[38] ), 
        .C(\B_DOUT_TEMPR97[38] ), .D(\B_DOUT_TEMPR98[38] ), .Y(
        OR4_610_Y));
    OR4 OR4_1403 (.A(\A_DOUT_TEMPR44[23] ), .B(\A_DOUT_TEMPR45[23] ), 
        .C(\A_DOUT_TEMPR46[23] ), .D(\A_DOUT_TEMPR47[23] ), .Y(
        OR4_1403_Y));
    OR4 OR4_1496 (.A(\B_DOUT_TEMPR107[34] ), .B(\B_DOUT_TEMPR108[34] ), 
        .C(\B_DOUT_TEMPR109[34] ), .D(\B_DOUT_TEMPR110[34] ), .Y(
        OR4_1496_Y));
    OR4 OR4_1058 (.A(\A_DOUT_TEMPR91[33] ), .B(\A_DOUT_TEMPR92[33] ), 
        .C(\A_DOUT_TEMPR93[33] ), .D(\A_DOUT_TEMPR94[33] ), .Y(
        OR4_1058_Y));
    OR4 OR4_808 (.A(\B_DOUT_TEMPR75[24] ), .B(\B_DOUT_TEMPR76[24] ), 
        .C(\B_DOUT_TEMPR77[24] ), .D(\B_DOUT_TEMPR78[24] ), .Y(
        OR4_808_Y));
    OR4 OR4_922 (.A(\A_DOUT_TEMPR12[20] ), .B(\A_DOUT_TEMPR13[20] ), 
        .C(\A_DOUT_TEMPR14[20] ), .D(\A_DOUT_TEMPR15[20] ), .Y(
        OR4_922_Y));
    OR4 OR4_601 (.A(\B_DOUT_TEMPR8[37] ), .B(\B_DOUT_TEMPR9[37] ), .C(
        \B_DOUT_TEMPR10[37] ), .D(\B_DOUT_TEMPR11[37] ), .Y(OR4_601_Y));
    OR4 OR4_647 (.A(\B_DOUT_TEMPR68[21] ), .B(\B_DOUT_TEMPR69[21] ), 
        .C(\B_DOUT_TEMPR70[21] ), .D(\B_DOUT_TEMPR71[21] ), .Y(
        OR4_647_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%50%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R50C1 (
        .A_DOUT({nc20820, nc20821, nc20822, nc20823, nc20824, nc20825, 
        nc20826, nc20827, nc20828, nc20829, nc20830, nc20831, nc20832, 
        nc20833, nc20834, \A_DOUT_TEMPR50[9] , \A_DOUT_TEMPR50[8] , 
        \A_DOUT_TEMPR50[7] , \A_DOUT_TEMPR50[6] , \A_DOUT_TEMPR50[5] })
        , .B_DOUT({nc20835, nc20836, nc20837, nc20838, nc20839, 
        nc20840, nc20841, nc20842, nc20843, nc20844, nc20845, nc20846, 
        nc20847, nc20848, nc20849, \B_DOUT_TEMPR50[9] , 
        \B_DOUT_TEMPR50[8] , \B_DOUT_TEMPR50[7] , \B_DOUT_TEMPR50[6] , 
        \B_DOUT_TEMPR50[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_125 (.A(OR4_668_Y), .B(OR4_1473_Y), .C(OR4_544_Y), .D(
        OR4_2892_Y), .Y(OR4_125_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%106%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R106C0 (
        .A_DOUT({nc20850, nc20851, nc20852, nc20853, nc20854, nc20855, 
        nc20856, nc20857, nc20858, nc20859, nc20860, nc20861, nc20862, 
        nc20863, nc20864, \A_DOUT_TEMPR106[4] , \A_DOUT_TEMPR106[3] , 
        \A_DOUT_TEMPR106[2] , \A_DOUT_TEMPR106[1] , 
        \A_DOUT_TEMPR106[0] }), .B_DOUT({nc20865, nc20866, nc20867, 
        nc20868, nc20869, nc20870, nc20871, nc20872, nc20873, nc20874, 
        nc20875, nc20876, nc20877, nc20878, nc20879, 
        \B_DOUT_TEMPR106[4] , \B_DOUT_TEMPR106[3] , 
        \B_DOUT_TEMPR106[2] , \B_DOUT_TEMPR106[1] , 
        \B_DOUT_TEMPR106[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[106][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1867 (.A(\A_DOUT_TEMPR111[28] ), .B(\A_DOUT_TEMPR112[28] ), 
        .C(\A_DOUT_TEMPR113[28] ), .D(\A_DOUT_TEMPR114[28] ), .Y(
        OR4_1867_Y));
    OR4 OR4_491 (.A(\B_DOUT_TEMPR12[25] ), .B(\B_DOUT_TEMPR13[25] ), 
        .C(\B_DOUT_TEMPR14[25] ), .D(\B_DOUT_TEMPR15[25] ), .Y(
        OR4_491_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%106%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R106C5 (
        .A_DOUT({nc20880, nc20881, nc20882, nc20883, nc20884, nc20885, 
        nc20886, nc20887, nc20888, nc20889, nc20890, nc20891, nc20892, 
        nc20893, nc20894, \A_DOUT_TEMPR106[29] , \A_DOUT_TEMPR106[28] , 
        \A_DOUT_TEMPR106[27] , \A_DOUT_TEMPR106[26] , 
        \A_DOUT_TEMPR106[25] }), .B_DOUT({nc20895, nc20896, nc20897, 
        nc20898, nc20899, nc20900, nc20901, nc20902, nc20903, nc20904, 
        nc20905, nc20906, nc20907, nc20908, nc20909, 
        \B_DOUT_TEMPR106[29] , \B_DOUT_TEMPR106[28] , 
        \B_DOUT_TEMPR106[27] , \B_DOUT_TEMPR106[26] , 
        \B_DOUT_TEMPR106[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[106][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_920 (.A(OR4_1025_Y), .B(OR4_2493_Y), .C(OR4_45_Y), .D(
        OR4_2913_Y), .Y(OR4_920_Y));
    OR4 OR4_2381 (.A(OR4_574_Y), .B(OR4_358_Y), .C(OR4_1075_Y), .D(
        OR4_1366_Y), .Y(OR4_2381_Y));
    OR4 OR4_1084 (.A(\A_DOUT_TEMPR40[11] ), .B(\A_DOUT_TEMPR41[11] ), 
        .C(\A_DOUT_TEMPR42[11] ), .D(\A_DOUT_TEMPR43[11] ), .Y(
        OR4_1084_Y));
    OR2 OR2_46 (.A(\B_DOUT_TEMPR72[25] ), .B(\B_DOUT_TEMPR73[25] ), .Y(
        OR2_46_Y));
    OR2 OR2_9 (.A(\A_DOUT_TEMPR72[1] ), .B(\A_DOUT_TEMPR73[1] ), .Y(
        OR2_9_Y));
    OR4 OR4_1086 (.A(\A_DOUT_TEMPR28[18] ), .B(\A_DOUT_TEMPR29[18] ), 
        .C(\A_DOUT_TEMPR30[18] ), .D(\A_DOUT_TEMPR31[18] ), .Y(
        OR4_1086_Y));
    OR4 OR4_859 (.A(OR4_991_Y), .B(OR4_1886_Y), .C(OR4_1529_Y), .D(
        OR4_0_Y), .Y(OR4_859_Y));
    OR4 OR4_1228 (.A(\B_DOUT_TEMPR83[27] ), .B(\B_DOUT_TEMPR84[27] ), 
        .C(\B_DOUT_TEMPR85[27] ), .D(\B_DOUT_TEMPR86[27] ), .Y(
        OR4_1228_Y));
    OR4 OR4_40 (.A(\A_DOUT_TEMPR40[18] ), .B(\A_DOUT_TEMPR41[18] ), .C(
        \A_DOUT_TEMPR42[18] ), .D(\A_DOUT_TEMPR43[18] ), .Y(OR4_40_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%5%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R5C6 (
        .A_DOUT({nc20910, nc20911, nc20912, nc20913, nc20914, nc20915, 
        nc20916, nc20917, nc20918, nc20919, nc20920, nc20921, nc20922, 
        nc20923, nc20924, \A_DOUT_TEMPR5[34] , \A_DOUT_TEMPR5[33] , 
        \A_DOUT_TEMPR5[32] , \A_DOUT_TEMPR5[31] , \A_DOUT_TEMPR5[30] })
        , .B_DOUT({nc20925, nc20926, nc20927, nc20928, nc20929, 
        nc20930, nc20931, nc20932, nc20933, nc20934, nc20935, nc20936, 
        nc20937, nc20938, nc20939, \B_DOUT_TEMPR5[34] , 
        \B_DOUT_TEMPR5[33] , \B_DOUT_TEMPR5[32] , \B_DOUT_TEMPR5[31] , 
        \B_DOUT_TEMPR5[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2881 (.A(OR4_2129_Y), .B(OR4_2485_Y), .C(OR4_1659_Y), .D(
        OR4_608_Y), .Y(OR4_2881_Y));
    OR4 OR4_1795 (.A(\B_DOUT_TEMPR111[35] ), .B(\B_DOUT_TEMPR112[35] ), 
        .C(\B_DOUT_TEMPR113[35] ), .D(\B_DOUT_TEMPR114[35] ), .Y(
        OR4_1795_Y));
    OR4 OR4_2174 (.A(\A_DOUT_TEMPR32[5] ), .B(\A_DOUT_TEMPR33[5] ), .C(
        \A_DOUT_TEMPR34[5] ), .D(\A_DOUT_TEMPR35[5] ), .Y(OR4_2174_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%33%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R33C3 (
        .A_DOUT({nc20940, nc20941, nc20942, nc20943, nc20944, nc20945, 
        nc20946, nc20947, nc20948, nc20949, nc20950, nc20951, nc20952, 
        nc20953, nc20954, \A_DOUT_TEMPR33[19] , \A_DOUT_TEMPR33[18] , 
        \A_DOUT_TEMPR33[17] , \A_DOUT_TEMPR33[16] , 
        \A_DOUT_TEMPR33[15] }), .B_DOUT({nc20955, nc20956, nc20957, 
        nc20958, nc20959, nc20960, nc20961, nc20962, nc20963, nc20964, 
        nc20965, nc20966, nc20967, nc20968, nc20969, 
        \B_DOUT_TEMPR33[19] , \B_DOUT_TEMPR33[18] , 
        \B_DOUT_TEMPR33[17] , \B_DOUT_TEMPR33[16] , 
        \B_DOUT_TEMPR33[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[33][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_404 (.A(\A_DOUT_TEMPR103[15] ), .B(\A_DOUT_TEMPR104[15] ), 
        .C(\A_DOUT_TEMPR105[15] ), .D(\A_DOUT_TEMPR106[15] ), .Y(
        OR4_404_Y));
    OR4 OR4_2951 (.A(\B_DOUT_TEMPR95[25] ), .B(\B_DOUT_TEMPR96[25] ), 
        .C(\B_DOUT_TEMPR97[25] ), .D(\B_DOUT_TEMPR98[25] ), .Y(
        OR4_2951_Y));
    OR4 OR4_251 (.A(\B_DOUT_TEMPR0[19] ), .B(\B_DOUT_TEMPR1[19] ), .C(
        \B_DOUT_TEMPR2[19] ), .D(\B_DOUT_TEMPR3[19] ), .Y(OR4_251_Y));
    OR4 OR4_851 (.A(OR4_1482_Y), .B(OR4_1786_Y), .C(OR4_1423_Y), .D(
        OR4_1806_Y), .Y(OR4_851_Y));
    OR4 OR4_2666 (.A(OR4_1990_Y), .B(OR4_2994_Y), .C(OR4_623_Y), .D(
        OR4_2270_Y), .Y(OR4_2666_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%35%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R35C3 (
        .A_DOUT({nc20970, nc20971, nc20972, nc20973, nc20974, nc20975, 
        nc20976, nc20977, nc20978, nc20979, nc20980, nc20981, nc20982, 
        nc20983, nc20984, \A_DOUT_TEMPR35[19] , \A_DOUT_TEMPR35[18] , 
        \A_DOUT_TEMPR35[17] , \A_DOUT_TEMPR35[16] , 
        \A_DOUT_TEMPR35[15] }), .B_DOUT({nc20985, nc20986, nc20987, 
        nc20988, nc20989, nc20990, nc20991, nc20992, nc20993, nc20994, 
        nc20995, nc20996, nc20997, nc20998, nc20999, 
        \B_DOUT_TEMPR35[19] , \B_DOUT_TEMPR35[18] , 
        \B_DOUT_TEMPR35[17] , \B_DOUT_TEMPR35[16] , 
        \B_DOUT_TEMPR35[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[35][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1213 (.A(OR4_1242_Y), .B(OR4_1023_Y), .C(OR4_2470_Y), .D(
        OR4_1027_Y), .Y(OR4_1213_Y));
    OR2 OR2_3 (.A(\B_DOUT_TEMPR72[17] ), .B(\B_DOUT_TEMPR73[17] ), .Y(
        OR2_3_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%111%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R111C2 (
        .A_DOUT({nc21000, nc21001, nc21002, nc21003, nc21004, nc21005, 
        nc21006, nc21007, nc21008, nc21009, nc21010, nc21011, nc21012, 
        nc21013, nc21014, \A_DOUT_TEMPR111[14] , \A_DOUT_TEMPR111[13] , 
        \A_DOUT_TEMPR111[12] , \A_DOUT_TEMPR111[11] , 
        \A_DOUT_TEMPR111[10] }), .B_DOUT({nc21015, nc21016, nc21017, 
        nc21018, nc21019, nc21020, nc21021, nc21022, nc21023, nc21024, 
        nc21025, nc21026, nc21027, nc21028, nc21029, 
        \B_DOUT_TEMPR111[14] , \B_DOUT_TEMPR111[13] , 
        \B_DOUT_TEMPR111[12] , \B_DOUT_TEMPR111[11] , 
        \B_DOUT_TEMPR111[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[111][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2160 (.A(\A_DOUT_TEMPR99[33] ), .B(\A_DOUT_TEMPR100[33] ), 
        .C(\A_DOUT_TEMPR101[33] ), .D(\A_DOUT_TEMPR102[33] ), .Y(
        OR4_2160_Y));
    OR4 OR4_1973 (.A(\B_DOUT_TEMPR60[38] ), .B(\B_DOUT_TEMPR61[38] ), 
        .C(\B_DOUT_TEMPR62[38] ), .D(\B_DOUT_TEMPR63[38] ), .Y(
        OR4_1973_Y));
    OR4 OR4_487 (.A(\B_DOUT_TEMPR83[34] ), .B(\B_DOUT_TEMPR84[34] ), 
        .C(\B_DOUT_TEMPR85[34] ), .D(\B_DOUT_TEMPR86[34] ), .Y(
        OR4_487_Y));
    OR4 OR4_65 (.A(\A_DOUT_TEMPR8[26] ), .B(\A_DOUT_TEMPR9[26] ), .C(
        \A_DOUT_TEMPR10[26] ), .D(\A_DOUT_TEMPR11[26] ), .Y(OR4_65_Y));
    OR4 OR4_1383 (.A(\A_DOUT_TEMPR28[6] ), .B(\A_DOUT_TEMPR29[6] ), .C(
        \A_DOUT_TEMPR30[6] ), .D(\A_DOUT_TEMPR31[6] ), .Y(OR4_1383_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%92%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R92C0 (
        .A_DOUT({nc21030, nc21031, nc21032, nc21033, nc21034, nc21035, 
        nc21036, nc21037, nc21038, nc21039, nc21040, nc21041, nc21042, 
        nc21043, nc21044, \A_DOUT_TEMPR92[4] , \A_DOUT_TEMPR92[3] , 
        \A_DOUT_TEMPR92[2] , \A_DOUT_TEMPR92[1] , \A_DOUT_TEMPR92[0] })
        , .B_DOUT({nc21045, nc21046, nc21047, nc21048, nc21049, 
        nc21050, nc21051, nc21052, nc21053, nc21054, nc21055, nc21056, 
        nc21057, nc21058, nc21059, \B_DOUT_TEMPR92[4] , 
        \B_DOUT_TEMPR92[3] , \B_DOUT_TEMPR92[2] , \B_DOUT_TEMPR92[1] , 
        \B_DOUT_TEMPR92[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[92][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1154 (.A(\A_DOUT_TEMPR60[38] ), .B(\A_DOUT_TEMPR61[38] ), 
        .C(\A_DOUT_TEMPR62[38] ), .D(\A_DOUT_TEMPR63[38] ), .Y(
        OR4_1154_Y));
    OR4 OR4_247 (.A(\A_DOUT_TEMPR107[31] ), .B(\A_DOUT_TEMPR108[31] ), 
        .C(\A_DOUT_TEMPR109[31] ), .D(\A_DOUT_TEMPR110[31] ), .Y(
        OR4_247_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%22%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R22C7 (
        .A_DOUT({nc21060, nc21061, nc21062, nc21063, nc21064, nc21065, 
        nc21066, nc21067, nc21068, nc21069, nc21070, nc21071, nc21072, 
        nc21073, nc21074, \A_DOUT_TEMPR22[39] , \A_DOUT_TEMPR22[38] , 
        \A_DOUT_TEMPR22[37] , \A_DOUT_TEMPR22[36] , 
        \A_DOUT_TEMPR22[35] }), .B_DOUT({nc21075, nc21076, nc21077, 
        nc21078, nc21079, nc21080, nc21081, nc21082, nc21083, nc21084, 
        nc21085, nc21086, nc21087, nc21088, nc21089, 
        \B_DOUT_TEMPR22[39] , \B_DOUT_TEMPR22[38] , 
        \B_DOUT_TEMPR22[37] , \B_DOUT_TEMPR22[36] , 
        \B_DOUT_TEMPR22[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%8%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R8C3 (
        .A_DOUT({nc21090, nc21091, nc21092, nc21093, nc21094, nc21095, 
        nc21096, nc21097, nc21098, nc21099, nc21100, nc21101, nc21102, 
        nc21103, nc21104, \A_DOUT_TEMPR8[19] , \A_DOUT_TEMPR8[18] , 
        \A_DOUT_TEMPR8[17] , \A_DOUT_TEMPR8[16] , \A_DOUT_TEMPR8[15] })
        , .B_DOUT({nc21105, nc21106, nc21107, nc21108, nc21109, 
        nc21110, nc21111, nc21112, nc21113, nc21114, nc21115, nc21116, 
        nc21117, nc21118, nc21119, \B_DOUT_TEMPR8[19] , 
        \B_DOUT_TEMPR8[18] , \B_DOUT_TEMPR8[17] , \B_DOUT_TEMPR8[16] , 
        \B_DOUT_TEMPR8[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_332 (.A(\B_DOUT_TEMPR75[5] ), .B(\B_DOUT_TEMPR76[5] ), .C(
        \B_DOUT_TEMPR77[5] ), .D(\B_DOUT_TEMPR78[5] ), .Y(OR4_332_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%91%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R91C6 (
        .A_DOUT({nc21120, nc21121, nc21122, nc21123, nc21124, nc21125, 
        nc21126, nc21127, nc21128, nc21129, nc21130, nc21131, nc21132, 
        nc21133, nc21134, \A_DOUT_TEMPR91[34] , \A_DOUT_TEMPR91[33] , 
        \A_DOUT_TEMPR91[32] , \A_DOUT_TEMPR91[31] , 
        \A_DOUT_TEMPR91[30] }), .B_DOUT({nc21135, nc21136, nc21137, 
        nc21138, nc21139, nc21140, nc21141, nc21142, nc21143, nc21144, 
        nc21145, nc21146, nc21147, nc21148, nc21149, 
        \B_DOUT_TEMPR91[34] , \B_DOUT_TEMPR91[33] , 
        \B_DOUT_TEMPR91[32] , \B_DOUT_TEMPR91[31] , 
        \B_DOUT_TEMPR91[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[91][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_874 (.A(\A_DOUT_TEMPR32[32] ), .B(\A_DOUT_TEMPR33[32] ), 
        .C(\A_DOUT_TEMPR34[32] ), .D(\A_DOUT_TEMPR35[32] ), .Y(
        OR4_874_Y));
    OR4 OR4_1371 (.A(\A_DOUT_TEMPR103[39] ), .B(\A_DOUT_TEMPR104[39] ), 
        .C(\A_DOUT_TEMPR105[39] ), .D(\A_DOUT_TEMPR106[39] ), .Y(
        OR4_1371_Y));
    OR4 OR4_2875 (.A(\A_DOUT_TEMPR64[7] ), .B(\A_DOUT_TEMPR65[7] ), .C(
        \A_DOUT_TEMPR66[7] ), .D(\A_DOUT_TEMPR67[7] ), .Y(OR4_2875_Y));
    OR4 OR4_2024 (.A(\B_DOUT_TEMPR24[9] ), .B(\B_DOUT_TEMPR25[9] ), .C(
        \B_DOUT_TEMPR26[9] ), .D(\B_DOUT_TEMPR27[9] ), .Y(OR4_2024_Y));
    OR4 \OR4_B_DOUT[37]  (.A(OR4_392_Y), .B(OR4_1381_Y), .C(OR4_1476_Y)
        , .D(OR4_1372_Y), .Y(B_DOUT[37]));
    OR4 OR4_2026 (.A(\A_DOUT_TEMPR28[13] ), .B(\A_DOUT_TEMPR29[13] ), 
        .C(\A_DOUT_TEMPR30[13] ), .D(\A_DOUT_TEMPR31[13] ), .Y(
        OR4_2026_Y));
    OR4 OR4_572 (.A(\A_DOUT_TEMPR12[38] ), .B(\A_DOUT_TEMPR13[38] ), 
        .C(\A_DOUT_TEMPR14[38] ), .D(\A_DOUT_TEMPR15[38] ), .Y(
        OR4_572_Y));
    OR4 OR4_1871 (.A(\A_DOUT_TEMPR4[2] ), .B(\A_DOUT_TEMPR5[2] ), .C(
        \A_DOUT_TEMPR6[2] ), .D(\A_DOUT_TEMPR7[2] ), .Y(OR4_1871_Y));
    OR4 OR4_2253 (.A(OR4_1796_Y), .B(OR4_2101_Y), .C(OR4_1724_Y), .D(
        OR4_2119_Y), .Y(OR4_2253_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%30%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R30C1 (
        .A_DOUT({nc21150, nc21151, nc21152, nc21153, nc21154, nc21155, 
        nc21156, nc21157, nc21158, nc21159, nc21160, nc21161, nc21162, 
        nc21163, nc21164, \A_DOUT_TEMPR30[9] , \A_DOUT_TEMPR30[8] , 
        \A_DOUT_TEMPR30[7] , \A_DOUT_TEMPR30[6] , \A_DOUT_TEMPR30[5] })
        , .B_DOUT({nc21165, nc21166, nc21167, nc21168, nc21169, 
        nc21170, nc21171, nc21172, nc21173, nc21174, nc21175, nc21176, 
        nc21177, nc21178, nc21179, \B_DOUT_TEMPR30[9] , 
        \B_DOUT_TEMPR30[8] , \B_DOUT_TEMPR30[7] , \B_DOUT_TEMPR30[6] , 
        \B_DOUT_TEMPR30[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_942 (.A(\B_DOUT_TEMPR56[25] ), .B(\B_DOUT_TEMPR57[25] ), 
        .C(\B_DOUT_TEMPR58[25] ), .D(\B_DOUT_TEMPR59[25] ), .Y(
        OR4_942_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%13%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R13C2 (
        .A_DOUT({nc21180, nc21181, nc21182, nc21183, nc21184, nc21185, 
        nc21186, nc21187, nc21188, nc21189, nc21190, nc21191, nc21192, 
        nc21193, nc21194, \A_DOUT_TEMPR13[14] , \A_DOUT_TEMPR13[13] , 
        \A_DOUT_TEMPR13[12] , \A_DOUT_TEMPR13[11] , 
        \A_DOUT_TEMPR13[10] }), .B_DOUT({nc21195, nc21196, nc21197, 
        nc21198, nc21199, nc21200, nc21201, nc21202, nc21203, nc21204, 
        nc21205, nc21206, nc21207, nc21208, nc21209, 
        \B_DOUT_TEMPR13[14] , \B_DOUT_TEMPR13[13] , 
        \B_DOUT_TEMPR13[12] , \B_DOUT_TEMPR13[11] , 
        \B_DOUT_TEMPR13[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%113%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R113C4 (
        .A_DOUT({nc21210, nc21211, nc21212, nc21213, nc21214, nc21215, 
        nc21216, nc21217, nc21218, nc21219, nc21220, nc21221, nc21222, 
        nc21223, nc21224, \A_DOUT_TEMPR113[24] , \A_DOUT_TEMPR113[23] , 
        \A_DOUT_TEMPR113[22] , \A_DOUT_TEMPR113[21] , 
        \A_DOUT_TEMPR113[20] }), .B_DOUT({nc21225, nc21226, nc21227, 
        nc21228, nc21229, nc21230, nc21231, nc21232, nc21233, nc21234, 
        nc21235, nc21236, nc21237, nc21238, nc21239, 
        \B_DOUT_TEMPR113[24] , \B_DOUT_TEMPR113[23] , 
        \B_DOUT_TEMPR113[22] , \B_DOUT_TEMPR113[21] , 
        \B_DOUT_TEMPR113[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[113][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_145 (.A(\A_DOUT_TEMPR115[29] ), .B(\A_DOUT_TEMPR116[29] ), 
        .C(\A_DOUT_TEMPR117[29] ), .D(\A_DOUT_TEMPR118[29] ), .Y(
        OR4_145_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%49%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R49C3 (
        .A_DOUT({nc21240, nc21241, nc21242, nc21243, nc21244, nc21245, 
        nc21246, nc21247, nc21248, nc21249, nc21250, nc21251, nc21252, 
        nc21253, nc21254, \A_DOUT_TEMPR49[19] , \A_DOUT_TEMPR49[18] , 
        \A_DOUT_TEMPR49[17] , \A_DOUT_TEMPR49[16] , 
        \A_DOUT_TEMPR49[15] }), .B_DOUT({nc21255, nc21256, nc21257, 
        nc21258, nc21259, nc21260, nc21261, nc21262, nc21263, nc21264, 
        nc21265, nc21266, nc21267, nc21268, nc21269, 
        \B_DOUT_TEMPR49[19] , \B_DOUT_TEMPR49[18] , 
        \B_DOUT_TEMPR49[17] , \B_DOUT_TEMPR49[16] , 
        \B_DOUT_TEMPR49[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[10]  (.A(OR4_439_Y), .B(OR4_2754_Y), .C(OR4_2934_Y)
        , .D(OR4_1256_Y), .Y(A_DOUT[10]));
    OR4 OR4_940 (.A(OR4_2772_Y), .B(OR4_2562_Y), .C(OR2_64_Y), .D(
        \A_DOUT_TEMPR74[31] ), .Y(OR4_940_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[4]  (.A(CFG3_4_Y), .B(CFG3_14_Y)
        , .Y(\BLKX2[4] ));
    OR4 OR4_1855 (.A(\B_DOUT_TEMPR64[23] ), .B(\B_DOUT_TEMPR65[23] ), 
        .C(\B_DOUT_TEMPR66[23] ), .D(\B_DOUT_TEMPR67[23] ), .Y(
        OR4_1855_Y));
    OR4 OR4_357 (.A(\A_DOUT_TEMPR40[12] ), .B(\A_DOUT_TEMPR41[12] ), 
        .C(\A_DOUT_TEMPR42[12] ), .D(\A_DOUT_TEMPR43[12] ), .Y(
        OR4_357_Y));
    OR4 OR4_2323 (.A(\A_DOUT_TEMPR107[32] ), .B(\A_DOUT_TEMPR108[32] ), 
        .C(\A_DOUT_TEMPR109[32] ), .D(\A_DOUT_TEMPR110[32] ), .Y(
        OR4_2323_Y));
    OR4 OR4_1941 (.A(\A_DOUT_TEMPR115[32] ), .B(\A_DOUT_TEMPR116[32] ), 
        .C(\A_DOUT_TEMPR117[32] ), .D(\A_DOUT_TEMPR118[32] ), .Y(
        OR4_1941_Y));
    OR4 OR4_858 (.A(\A_DOUT_TEMPR56[16] ), .B(\A_DOUT_TEMPR57[16] ), 
        .C(\A_DOUT_TEMPR58[16] ), .D(\A_DOUT_TEMPR59[16] ), .Y(
        OR4_858_Y));
    OR4 \OR4_B_DOUT[25]  (.A(OR4_1825_Y), .B(OR4_2064_Y), .C(
        OR4_2873_Y), .D(OR4_636_Y), .Y(B_DOUT[25]));
    OR4 OR4_2249 (.A(OR4_1555_Y), .B(OR4_1018_Y), .C(OR4_1620_Y), .D(
        OR4_814_Y), .Y(OR4_2249_Y));
    OR4 OR4_651 (.A(\B_DOUT_TEMPR4[36] ), .B(\B_DOUT_TEMPR5[36] ), .C(
        \B_DOUT_TEMPR6[36] ), .D(\B_DOUT_TEMPR7[36] ), .Y(OR4_651_Y));
    OR4 OR4_1206 (.A(\A_DOUT_TEMPR0[30] ), .B(\A_DOUT_TEMPR1[30] ), .C(
        \A_DOUT_TEMPR2[30] ), .D(\A_DOUT_TEMPR3[30] ), .Y(OR4_1206_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%1%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R1C7 (
        .A_DOUT({nc21270, nc21271, nc21272, nc21273, nc21274, nc21275, 
        nc21276, nc21277, nc21278, nc21279, nc21280, nc21281, nc21282, 
        nc21283, nc21284, \A_DOUT_TEMPR1[39] , \A_DOUT_TEMPR1[38] , 
        \A_DOUT_TEMPR1[37] , \A_DOUT_TEMPR1[36] , \A_DOUT_TEMPR1[35] })
        , .B_DOUT({nc21285, nc21286, nc21287, nc21288, nc21289, 
        nc21290, nc21291, nc21292, nc21293, nc21294, nc21295, nc21296, 
        nc21297, nc21298, nc21299, \B_DOUT_TEMPR1[39] , 
        \B_DOUT_TEMPR1[38] , \B_DOUT_TEMPR1[37] , \B_DOUT_TEMPR1[36] , 
        \B_DOUT_TEMPR1[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_535 (.A(\B_DOUT_TEMPR95[28] ), .B(\B_DOUT_TEMPR96[28] ), 
        .C(\B_DOUT_TEMPR97[28] ), .D(\B_DOUT_TEMPR98[28] ), .Y(
        OR4_535_Y));
    OR4 OR4_2635 (.A(\B_DOUT_TEMPR64[32] ), .B(\B_DOUT_TEMPR65[32] ), 
        .C(\B_DOUT_TEMPR66[32] ), .D(\B_DOUT_TEMPR67[32] ), .Y(
        OR4_2635_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%98%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R98C2 (
        .A_DOUT({nc21300, nc21301, nc21302, nc21303, nc21304, nc21305, 
        nc21306, nc21307, nc21308, nc21309, nc21310, nc21311, nc21312, 
        nc21313, nc21314, \A_DOUT_TEMPR98[14] , \A_DOUT_TEMPR98[13] , 
        \A_DOUT_TEMPR98[12] , \A_DOUT_TEMPR98[11] , 
        \A_DOUT_TEMPR98[10] }), .B_DOUT({nc21315, nc21316, nc21317, 
        nc21318, nc21319, nc21320, nc21321, nc21322, nc21323, nc21324, 
        nc21325, nc21326, nc21327, nc21328, nc21329, 
        \B_DOUT_TEMPR98[14] , \B_DOUT_TEMPR98[13] , 
        \B_DOUT_TEMPR98[12] , \B_DOUT_TEMPR98[11] , 
        \B_DOUT_TEMPR98[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[98][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%47%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R47C3 (
        .A_DOUT({nc21330, nc21331, nc21332, nc21333, nc21334, nc21335, 
        nc21336, nc21337, nc21338, nc21339, nc21340, nc21341, nc21342, 
        nc21343, nc21344, \A_DOUT_TEMPR47[19] , \A_DOUT_TEMPR47[18] , 
        \A_DOUT_TEMPR47[17] , \A_DOUT_TEMPR47[16] , 
        \A_DOUT_TEMPR47[15] }), .B_DOUT({nc21345, nc21346, nc21347, 
        nc21348, nc21349, nc21350, nc21351, nc21352, nc21353, nc21354, 
        nc21355, nc21356, nc21357, nc21358, nc21359, 
        \B_DOUT_TEMPR47[19] , \B_DOUT_TEMPR47[18] , 
        \B_DOUT_TEMPR47[17] , \B_DOUT_TEMPR47[16] , 
        \B_DOUT_TEMPR47[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%50%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R50C7 (
        .A_DOUT({nc21360, nc21361, nc21362, nc21363, nc21364, nc21365, 
        nc21366, nc21367, nc21368, nc21369, nc21370, nc21371, nc21372, 
        nc21373, nc21374, \A_DOUT_TEMPR50[39] , \A_DOUT_TEMPR50[38] , 
        \A_DOUT_TEMPR50[37] , \A_DOUT_TEMPR50[36] , 
        \A_DOUT_TEMPR50[35] }), .B_DOUT({nc21375, nc21376, nc21377, 
        nc21378, nc21379, nc21380, nc21381, nc21382, nc21383, nc21384, 
        nc21385, nc21386, nc21387, nc21388, nc21389, 
        \B_DOUT_TEMPR50[39] , \B_DOUT_TEMPR50[38] , 
        \B_DOUT_TEMPR50[37] , \B_DOUT_TEMPR50[36] , 
        \B_DOUT_TEMPR50[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2997 (.A(OR4_1671_Y), .B(OR4_1032_Y), .C(OR2_76_Y), .D(
        \B_DOUT_TEMPR74[1] ), .Y(OR4_2997_Y));
    OR4 OR4_45 (.A(\A_DOUT_TEMPR24[31] ), .B(\A_DOUT_TEMPR25[31] ), .C(
        \A_DOUT_TEMPR26[31] ), .D(\A_DOUT_TEMPR27[31] ), .Y(OR4_45_Y));
    OR4 OR4_1635 (.A(OR4_2585_Y), .B(OR4_1355_Y), .C(OR4_990_Y), .D(
        OR4_2406_Y), .Y(OR4_1635_Y));
    OR4 OR4_804 (.A(\A_DOUT_TEMPR87[37] ), .B(\A_DOUT_TEMPR88[37] ), 
        .C(\A_DOUT_TEMPR89[37] ), .D(\A_DOUT_TEMPR90[37] ), .Y(
        OR4_804_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%19%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R19C4 (
        .A_DOUT({nc21390, nc21391, nc21392, nc21393, nc21394, nc21395, 
        nc21396, nc21397, nc21398, nc21399, nc21400, nc21401, nc21402, 
        nc21403, nc21404, \A_DOUT_TEMPR19[24] , \A_DOUT_TEMPR19[23] , 
        \A_DOUT_TEMPR19[22] , \A_DOUT_TEMPR19[21] , 
        \A_DOUT_TEMPR19[20] }), .B_DOUT({nc21405, nc21406, nc21407, 
        nc21408, nc21409, nc21410, nc21411, nc21412, nc21413, nc21414, 
        nc21415, nc21416, nc21417, nc21418, nc21419, 
        \B_DOUT_TEMPR19[24] , \B_DOUT_TEMPR19[23] , 
        \B_DOUT_TEMPR19[22] , \B_DOUT_TEMPR19[21] , 
        \B_DOUT_TEMPR19[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[19][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_260 (.A(\B_DOUT_TEMPR64[6] ), .B(\B_DOUT_TEMPR65[6] ), .C(
        \B_DOUT_TEMPR66[6] ), .D(\B_DOUT_TEMPR67[6] ), .Y(OR4_260_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%74%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R74C0 (
        .A_DOUT({nc21420, nc21421, nc21422, nc21423, nc21424, nc21425, 
        nc21426, nc21427, nc21428, nc21429, nc21430, nc21431, nc21432, 
        nc21433, nc21434, \A_DOUT_TEMPR74[4] , \A_DOUT_TEMPR74[3] , 
        \A_DOUT_TEMPR74[2] , \A_DOUT_TEMPR74[1] , \A_DOUT_TEMPR74[0] })
        , .B_DOUT({nc21435, nc21436, nc21437, nc21438, nc21439, 
        nc21440, nc21441, nc21442, nc21443, nc21444, nc21445, nc21446, 
        nc21447, nc21448, nc21449, \B_DOUT_TEMPR74[4] , 
        \B_DOUT_TEMPR74[3] , \B_DOUT_TEMPR74[2] , \B_DOUT_TEMPR74[1] , 
        \B_DOUT_TEMPR74[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[74][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1596 (.A(\B_DOUT_TEMPR8[22] ), .B(\B_DOUT_TEMPR9[22] ), .C(
        \B_DOUT_TEMPR10[22] ), .D(\B_DOUT_TEMPR11[22] ), .Y(OR4_1596_Y)
        );
    OR4 OR4_502 (.A(\A_DOUT_TEMPR0[17] ), .B(\A_DOUT_TEMPR1[17] ), .C(
        \A_DOUT_TEMPR2[17] ), .D(\A_DOUT_TEMPR3[17] ), .Y(OR4_502_Y));
    OR4 OR4_2963 (.A(\B_DOUT_TEMPR44[15] ), .B(\B_DOUT_TEMPR45[15] ), 
        .C(\B_DOUT_TEMPR46[15] ), .D(\B_DOUT_TEMPR47[15] ), .Y(
        OR4_2963_Y));
    OR4 OR4_454 (.A(OR4_2875_Y), .B(OR4_1258_Y), .C(OR2_25_Y), .D(
        \A_DOUT_TEMPR74[7] ), .Y(OR4_454_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%81%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R81C0 (
        .A_DOUT({nc21450, nc21451, nc21452, nc21453, nc21454, nc21455, 
        nc21456, nc21457, nc21458, nc21459, nc21460, nc21461, nc21462, 
        nc21463, nc21464, \A_DOUT_TEMPR81[4] , \A_DOUT_TEMPR81[3] , 
        \A_DOUT_TEMPR81[2] , \A_DOUT_TEMPR81[1] , \A_DOUT_TEMPR81[0] })
        , .B_DOUT({nc21465, nc21466, nc21467, nc21468, nc21469, 
        nc21470, nc21471, nc21472, nc21473, nc21474, nc21475, nc21476, 
        nc21477, nc21478, nc21479, \B_DOUT_TEMPR81[4] , 
        \B_DOUT_TEMPR81[3] , \B_DOUT_TEMPR81[2] , \B_DOUT_TEMPR81[1] , 
        \B_DOUT_TEMPR81[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[81][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_660 (.A(OR4_1938_Y), .B(OR4_2778_Y), .C(OR4_1807_Y), .D(
        OR4_997_Y), .Y(OR4_660_Y));
    OR4 OR4_1797 (.A(\A_DOUT_TEMPR8[12] ), .B(\A_DOUT_TEMPR9[12] ), .C(
        \A_DOUT_TEMPR10[12] ), .D(\A_DOUT_TEMPR11[12] ), .Y(OR4_1797_Y)
        );
    OR4 OR4_3030 (.A(\A_DOUT_TEMPR103[38] ), .B(\A_DOUT_TEMPR104[38] ), 
        .C(\A_DOUT_TEMPR105[38] ), .D(\A_DOUT_TEMPR106[38] ), .Y(
        OR4_3030_Y));
    OR4 OR4_899 (.A(OR4_2668_Y), .B(OR4_807_Y), .C(OR4_1851_Y), .D(
        OR4_2134_Y), .Y(OR4_899_Y));
    OR4 OR4_1591 (.A(\B_DOUT_TEMPR115[33] ), .B(\B_DOUT_TEMPR116[33] ), 
        .C(\B_DOUT_TEMPR117[33] ), .D(\B_DOUT_TEMPR118[33] ), .Y(
        OR4_1591_Y));
    OR4 OR4_1243 (.A(\B_DOUT_TEMPR28[30] ), .B(\B_DOUT_TEMPR29[30] ), 
        .C(\B_DOUT_TEMPR30[30] ), .D(\B_DOUT_TEMPR31[30] ), .Y(
        OR4_1243_Y));
    OR4 OR4_2637 (.A(\B_DOUT_TEMPR68[6] ), .B(\B_DOUT_TEMPR69[6] ), .C(
        \B_DOUT_TEMPR70[6] ), .D(\B_DOUT_TEMPR71[6] ), .Y(OR4_2637_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%98%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R98C3 (
        .A_DOUT({nc21480, nc21481, nc21482, nc21483, nc21484, nc21485, 
        nc21486, nc21487, nc21488, nc21489, nc21490, nc21491, nc21492, 
        nc21493, nc21494, \A_DOUT_TEMPR98[19] , \A_DOUT_TEMPR98[18] , 
        \A_DOUT_TEMPR98[17] , \A_DOUT_TEMPR98[16] , 
        \A_DOUT_TEMPR98[15] }), .B_DOUT({nc21495, nc21496, nc21497, 
        nc21498, nc21499, nc21500, nc21501, nc21502, nc21503, nc21504, 
        nc21505, nc21506, nc21507, nc21508, nc21509, 
        \B_DOUT_TEMPR98[19] , \B_DOUT_TEMPR98[18] , 
        \B_DOUT_TEMPR98[17] , \B_DOUT_TEMPR98[16] , 
        \B_DOUT_TEMPR98[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[98][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_291 (.A(\A_DOUT_TEMPR83[29] ), .B(\A_DOUT_TEMPR84[29] ), 
        .C(\A_DOUT_TEMPR85[29] ), .D(\A_DOUT_TEMPR86[29] ), .Y(
        OR4_291_Y));
    OR4 OR4_2210 (.A(OR4_2112_Y), .B(OR4_2413_Y), .C(OR4_2052_Y), .D(
        OR4_2428_Y), .Y(OR4_2210_Y));
    OR4 OR4_891 (.A(OR4_854_Y), .B(OR4_1754_Y), .C(OR4_1410_Y), .D(
        OR4_2931_Y), .Y(OR4_891_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%76%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R76C7 (
        .A_DOUT({nc21510, nc21511, nc21512, nc21513, nc21514, nc21515, 
        nc21516, nc21517, nc21518, nc21519, nc21520, nc21521, nc21522, 
        nc21523, nc21524, \A_DOUT_TEMPR76[39] , \A_DOUT_TEMPR76[38] , 
        \A_DOUT_TEMPR76[37] , \A_DOUT_TEMPR76[36] , 
        \A_DOUT_TEMPR76[35] }), .B_DOUT({nc21525, nc21526, nc21527, 
        nc21528, nc21529, nc21530, nc21531, nc21532, nc21533, nc21534, 
        nc21535, nc21536, nc21537, nc21538, nc21539, 
        \B_DOUT_TEMPR76[39] , \B_DOUT_TEMPR76[38] , 
        \B_DOUT_TEMPR76[37] , \B_DOUT_TEMPR76[36] , 
        \B_DOUT_TEMPR76[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[76][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%8%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R8C5 (
        .A_DOUT({nc21540, nc21541, nc21542, nc21543, nc21544, nc21545, 
        nc21546, nc21547, nc21548, nc21549, nc21550, nc21551, nc21552, 
        nc21553, nc21554, \A_DOUT_TEMPR8[29] , \A_DOUT_TEMPR8[28] , 
        \A_DOUT_TEMPR8[27] , \A_DOUT_TEMPR8[26] , \A_DOUT_TEMPR8[25] })
        , .B_DOUT({nc21555, nc21556, nc21557, nc21558, nc21559, 
        nc21560, nc21561, nc21562, nc21563, nc21564, nc21565, nc21566, 
        nc21567, nc21568, nc21569, \B_DOUT_TEMPR8[29] , 
        \B_DOUT_TEMPR8[28] , \B_DOUT_TEMPR8[27] , \B_DOUT_TEMPR8[26] , 
        \B_DOUT_TEMPR8[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1637 (.A(\B_DOUT_TEMPR87[3] ), .B(\B_DOUT_TEMPR88[3] ), .C(
        \B_DOUT_TEMPR89[3] ), .D(\B_DOUT_TEMPR90[3] ), .Y(OR4_1637_Y));
    OR4 OR4_2987 (.A(\B_DOUT_TEMPR87[17] ), .B(\B_DOUT_TEMPR88[17] ), 
        .C(\B_DOUT_TEMPR89[17] ), .D(\B_DOUT_TEMPR90[17] ), .Y(
        OR4_2987_Y));
    OR4 OR4_2361 (.A(\B_DOUT_TEMPR16[30] ), .B(\B_DOUT_TEMPR17[30] ), 
        .C(\B_DOUT_TEMPR18[30] ), .D(\B_DOUT_TEMPR19[30] ), .Y(
        OR4_2361_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%94%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R94C1 (
        .A_DOUT({nc21570, nc21571, nc21572, nc21573, nc21574, nc21575, 
        nc21576, nc21577, nc21578, nc21579, nc21580, nc21581, nc21582, 
        nc21583, nc21584, \A_DOUT_TEMPR94[9] , \A_DOUT_TEMPR94[8] , 
        \A_DOUT_TEMPR94[7] , \A_DOUT_TEMPR94[6] , \A_DOUT_TEMPR94[5] })
        , .B_DOUT({nc21585, nc21586, nc21587, nc21588, nc21589, 
        nc21590, nc21591, nc21592, nc21593, nc21594, nc21595, nc21596, 
        nc21597, nc21598, nc21599, \B_DOUT_TEMPR94[9] , 
        \B_DOUT_TEMPR94[8] , \B_DOUT_TEMPR94[7] , \B_DOUT_TEMPR94[6] , 
        \B_DOUT_TEMPR94[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[94][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_69 (.A(\B_DOUT_TEMPR75[37] ), .B(\B_DOUT_TEMPR76[37] ), .C(
        \B_DOUT_TEMPR77[37] ), .D(\B_DOUT_TEMPR78[37] ), .Y(OR4_69_Y));
    OR4 OR4_2890 (.A(\A_DOUT_TEMPR28[21] ), .B(\A_DOUT_TEMPR29[21] ), 
        .C(\A_DOUT_TEMPR30[21] ), .D(\A_DOUT_TEMPR31[21] ), .Y(
        OR4_2890_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%90%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R90C4 (
        .A_DOUT({nc21600, nc21601, nc21602, nc21603, nc21604, nc21605, 
        nc21606, nc21607, nc21608, nc21609, nc21610, nc21611, nc21612, 
        nc21613, nc21614, \A_DOUT_TEMPR90[24] , \A_DOUT_TEMPR90[23] , 
        \A_DOUT_TEMPR90[22] , \A_DOUT_TEMPR90[21] , 
        \A_DOUT_TEMPR90[20] }), .B_DOUT({nc21615, nc21616, nc21617, 
        nc21618, nc21619, nc21620, nc21621, nc21622, nc21623, nc21624, 
        nc21625, nc21626, nc21627, nc21628, nc21629, 
        \B_DOUT_TEMPR90[24] , \B_DOUT_TEMPR90[23] , 
        \B_DOUT_TEMPR90[22] , \B_DOUT_TEMPR90[21] , 
        \B_DOUT_TEMPR90[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[90][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%63%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R63C3 (
        .A_DOUT({nc21630, nc21631, nc21632, nc21633, nc21634, nc21635, 
        nc21636, nc21637, nc21638, nc21639, nc21640, nc21641, nc21642, 
        nc21643, nc21644, \A_DOUT_TEMPR63[19] , \A_DOUT_TEMPR63[18] , 
        \A_DOUT_TEMPR63[17] , \A_DOUT_TEMPR63[16] , 
        \A_DOUT_TEMPR63[15] }), .B_DOUT({nc21645, nc21646, nc21647, 
        nc21648, nc21649, nc21650, nc21651, nc21652, nc21653, nc21654, 
        nc21655, nc21656, nc21657, nc21658, nc21659, 
        \B_DOUT_TEMPR63[19] , \B_DOUT_TEMPR63[18] , 
        \B_DOUT_TEMPR63[17] , \B_DOUT_TEMPR63[16] , 
        \B_DOUT_TEMPR63[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[63][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%77%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R77C6 (
        .A_DOUT({nc21660, nc21661, nc21662, nc21663, nc21664, nc21665, 
        nc21666, nc21667, nc21668, nc21669, nc21670, nc21671, nc21672, 
        nc21673, nc21674, \A_DOUT_TEMPR77[34] , \A_DOUT_TEMPR77[33] , 
        \A_DOUT_TEMPR77[32] , \A_DOUT_TEMPR77[31] , 
        \A_DOUT_TEMPR77[30] }), .B_DOUT({nc21675, nc21676, nc21677, 
        nc21678, nc21679, nc21680, nc21681, nc21682, nc21683, nc21684, 
        nc21685, nc21686, nc21687, nc21688, nc21689, 
        \B_DOUT_TEMPR77[34] , \B_DOUT_TEMPR77[33] , 
        \B_DOUT_TEMPR77[32] , \B_DOUT_TEMPR77[31] , 
        \B_DOUT_TEMPR77[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[77][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1806 (.A(\A_DOUT_TEMPR60[24] ), .B(\A_DOUT_TEMPR61[24] ), 
        .C(\A_DOUT_TEMPR62[24] ), .D(\A_DOUT_TEMPR63[24] ), .Y(
        OR4_1806_Y));
    OR4 OR4_2861 (.A(\B_DOUT_TEMPR83[16] ), .B(\B_DOUT_TEMPR84[16] ), 
        .C(\B_DOUT_TEMPR85[16] ), .D(\B_DOUT_TEMPR86[16] ), .Y(
        OR4_2861_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%65%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R65C3 (
        .A_DOUT({nc21690, nc21691, nc21692, nc21693, nc21694, nc21695, 
        nc21696, nc21697, nc21698, nc21699, nc21700, nc21701, nc21702, 
        nc21703, nc21704, \A_DOUT_TEMPR65[19] , \A_DOUT_TEMPR65[18] , 
        \A_DOUT_TEMPR65[17] , \A_DOUT_TEMPR65[16] , 
        \A_DOUT_TEMPR65[15] }), .B_DOUT({nc21705, nc21706, nc21707, 
        nc21708, nc21709, nc21710, nc21711, nc21712, nc21713, nc21714, 
        nc21715, nc21716, nc21717, nc21718, nc21719, 
        \B_DOUT_TEMPR65[19] , \B_DOUT_TEMPR65[18] , 
        \B_DOUT_TEMPR65[17] , \B_DOUT_TEMPR65[16] , 
        \B_DOUT_TEMPR65[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[65][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2503 (.A(\A_DOUT_TEMPR40[21] ), .B(\A_DOUT_TEMPR41[21] ), 
        .C(\A_DOUT_TEMPR42[21] ), .D(\A_DOUT_TEMPR43[21] ), .Y(
        OR4_2503_Y));
    OR4 OR4_2894 (.A(\B_DOUT_TEMPR64[21] ), .B(\B_DOUT_TEMPR65[21] ), 
        .C(\B_DOUT_TEMPR66[21] ), .D(\B_DOUT_TEMPR67[21] ), .Y(
        OR4_2894_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%107%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R107C2 (
        .A_DOUT({nc21720, nc21721, nc21722, nc21723, nc21724, nc21725, 
        nc21726, nc21727, nc21728, nc21729, nc21730, nc21731, nc21732, 
        nc21733, nc21734, \A_DOUT_TEMPR107[14] , \A_DOUT_TEMPR107[13] , 
        \A_DOUT_TEMPR107[12] , \A_DOUT_TEMPR107[11] , 
        \A_DOUT_TEMPR107[10] }), .B_DOUT({nc21735, nc21736, nc21737, 
        nc21738, nc21739, nc21740, nc21741, nc21742, nc21743, nc21744, 
        nc21745, nc21746, nc21747, nc21748, nc21749, 
        \B_DOUT_TEMPR107[14] , \B_DOUT_TEMPR107[13] , 
        \B_DOUT_TEMPR107[12] , \B_DOUT_TEMPR107[11] , 
        \B_DOUT_TEMPR107[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[107][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%111%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R111C6 (
        .A_DOUT({nc21750, nc21751, nc21752, nc21753, nc21754, nc21755, 
        nc21756, nc21757, nc21758, nc21759, nc21760, nc21761, nc21762, 
        nc21763, nc21764, \A_DOUT_TEMPR111[34] , \A_DOUT_TEMPR111[33] , 
        \A_DOUT_TEMPR111[32] , \A_DOUT_TEMPR111[31] , 
        \A_DOUT_TEMPR111[30] }), .B_DOUT({nc21765, nc21766, nc21767, 
        nc21768, nc21769, nc21770, nc21771, nc21772, nc21773, nc21774, 
        nc21775, nc21776, nc21777, nc21778, nc21779, 
        \B_DOUT_TEMPR111[34] , \B_DOUT_TEMPR111[33] , 
        \B_DOUT_TEMPR111[32] , \B_DOUT_TEMPR111[31] , 
        \B_DOUT_TEMPR111[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[111][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%72%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R72C4 (
        .A_DOUT({nc21780, nc21781, nc21782, nc21783, nc21784, nc21785, 
        nc21786, nc21787, nc21788, nc21789, nc21790, nc21791, nc21792, 
        nc21793, nc21794, \A_DOUT_TEMPR72[24] , \A_DOUT_TEMPR72[23] , 
        \A_DOUT_TEMPR72[22] , \A_DOUT_TEMPR72[21] , 
        \A_DOUT_TEMPR72[20] }), .B_DOUT({nc21795, nc21796, nc21797, 
        nc21798, nc21799, nc21800, nc21801, nc21802, nc21803, nc21804, 
        nc21805, nc21806, nc21807, nc21808, nc21809, 
        \B_DOUT_TEMPR72[24] , \B_DOUT_TEMPR72[23] , 
        \B_DOUT_TEMPR72[22] , \B_DOUT_TEMPR72[21] , 
        \B_DOUT_TEMPR72[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[72][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2103 (.A(\A_DOUT_TEMPR32[18] ), .B(\A_DOUT_TEMPR33[18] ), 
        .C(\A_DOUT_TEMPR34[18] ), .D(\A_DOUT_TEMPR35[18] ), .Y(
        OR4_2103_Y));
    OR4 OR4_2316 (.A(OR4_91_Y), .B(OR4_2105_Y), .C(OR4_2766_Y), .D(
        OR4_1933_Y), .Y(OR4_2316_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%111%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R111C7 (
        .A_DOUT({nc21810, nc21811, nc21812, nc21813, nc21814, nc21815, 
        nc21816, nc21817, nc21818, nc21819, nc21820, nc21821, nc21822, 
        nc21823, nc21824, \A_DOUT_TEMPR111[39] , \A_DOUT_TEMPR111[38] , 
        \A_DOUT_TEMPR111[37] , \A_DOUT_TEMPR111[36] , 
        \A_DOUT_TEMPR111[35] }), .B_DOUT({nc21825, nc21826, nc21827, 
        nc21828, nc21829, nc21830, nc21831, nc21832, nc21833, nc21834, 
        nc21835, nc21836, nc21837, nc21838, nc21839, 
        \B_DOUT_TEMPR111[39] , \B_DOUT_TEMPR111[38] , 
        \B_DOUT_TEMPR111[37] , \B_DOUT_TEMPR111[36] , 
        \B_DOUT_TEMPR111[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[111][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%3%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R3C4 (
        .A_DOUT({nc21840, nc21841, nc21842, nc21843, nc21844, nc21845, 
        nc21846, nc21847, nc21848, nc21849, nc21850, nc21851, nc21852, 
        nc21853, nc21854, \A_DOUT_TEMPR3[24] , \A_DOUT_TEMPR3[23] , 
        \A_DOUT_TEMPR3[22] , \A_DOUT_TEMPR3[21] , \A_DOUT_TEMPR3[20] })
        , .B_DOUT({nc21855, nc21856, nc21857, nc21858, nc21859, 
        nc21860, nc21861, nc21862, nc21863, nc21864, nc21865, nc21866, 
        nc21867, nc21868, nc21869, \B_DOUT_TEMPR3[24] , 
        \B_DOUT_TEMPR3[23] , \B_DOUT_TEMPR3[22] , \B_DOUT_TEMPR3[21] , 
        \B_DOUT_TEMPR3[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%30%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R30C7 (
        .A_DOUT({nc21870, nc21871, nc21872, nc21873, nc21874, nc21875, 
        nc21876, nc21877, nc21878, nc21879, nc21880, nc21881, nc21882, 
        nc21883, nc21884, \A_DOUT_TEMPR30[39] , \A_DOUT_TEMPR30[38] , 
        \A_DOUT_TEMPR30[37] , \A_DOUT_TEMPR30[36] , 
        \A_DOUT_TEMPR30[35] }), .B_DOUT({nc21885, nc21886, nc21887, 
        nc21888, nc21889, nc21890, nc21891, nc21892, nc21893, nc21894, 
        nc21895, nc21896, nc21897, nc21898, nc21899, 
        \B_DOUT_TEMPR30[39] , \B_DOUT_TEMPR30[38] , 
        \B_DOUT_TEMPR30[37] , \B_DOUT_TEMPR30[36] , 
        \B_DOUT_TEMPR30[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2002 (.A(\B_DOUT_TEMPR12[15] ), .B(\B_DOUT_TEMPR13[15] ), 
        .C(\B_DOUT_TEMPR14[15] ), .D(\B_DOUT_TEMPR15[15] ), .Y(
        OR4_2002_Y));
    OR4 OR4_2880 (.A(OR4_591_Y), .B(OR4_1579_Y), .C(OR4_2237_Y), .D(
        OR4_900_Y), .Y(OR4_2880_Y));
    OR4 OR4_1522 (.A(\B_DOUT_TEMPR48[30] ), .B(\B_DOUT_TEMPR49[30] ), 
        .C(\B_DOUT_TEMPR50[30] ), .D(\B_DOUT_TEMPR51[30] ), .Y(
        OR4_1522_Y));
    OR4 OR4_2678 (.A(\B_DOUT_TEMPR24[22] ), .B(\B_DOUT_TEMPR25[22] ), 
        .C(\B_DOUT_TEMPR26[22] ), .D(\B_DOUT_TEMPR27[22] ), .Y(
        OR4_2678_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%52%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R52C0 (
        .A_DOUT({nc21900, nc21901, nc21902, nc21903, nc21904, nc21905, 
        nc21906, nc21907, nc21908, nc21909, nc21910, nc21911, nc21912, 
        nc21913, nc21914, \A_DOUT_TEMPR52[4] , \A_DOUT_TEMPR52[3] , 
        \A_DOUT_TEMPR52[2] , \A_DOUT_TEMPR52[1] , \A_DOUT_TEMPR52[0] })
        , .B_DOUT({nc21915, nc21916, nc21917, nc21918, nc21919, 
        nc21920, nc21921, nc21922, nc21923, nc21924, nc21925, nc21926, 
        nc21927, nc21928, nc21929, \B_DOUT_TEMPR52[4] , 
        \B_DOUT_TEMPR52[3] , \B_DOUT_TEMPR52[2] , \B_DOUT_TEMPR52[1] , 
        \B_DOUT_TEMPR52[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[52][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1977 (.A(\B_DOUT_TEMPR95[15] ), .B(\B_DOUT_TEMPR96[15] ), 
        .C(\B_DOUT_TEMPR97[15] ), .D(\B_DOUT_TEMPR98[15] ), .Y(
        OR4_1977_Y));
    OR4 OR4_2884 (.A(\A_DOUT_TEMPR99[30] ), .B(\A_DOUT_TEMPR100[30] ), 
        .C(\A_DOUT_TEMPR101[30] ), .D(\A_DOUT_TEMPR102[30] ), .Y(
        OR4_2884_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%60%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R60C1 (
        .A_DOUT({nc21930, nc21931, nc21932, nc21933, nc21934, nc21935, 
        nc21936, nc21937, nc21938, nc21939, nc21940, nc21941, nc21942, 
        nc21943, nc21944, \A_DOUT_TEMPR60[9] , \A_DOUT_TEMPR60[8] , 
        \A_DOUT_TEMPR60[7] , \A_DOUT_TEMPR60[6] , \A_DOUT_TEMPR60[5] })
        , .B_DOUT({nc21945, nc21946, nc21947, nc21948, nc21949, 
        nc21950, nc21951, nc21952, nc21953, nc21954, nc21955, nc21956, 
        nc21957, nc21958, nc21959, \B_DOUT_TEMPR60[9] , 
        \B_DOUT_TEMPR60[8] , \B_DOUT_TEMPR60[7] , \B_DOUT_TEMPR60[6] , 
        \B_DOUT_TEMPR60[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[60][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1700 (.A(\A_DOUT_TEMPR99[21] ), .B(\A_DOUT_TEMPR100[21] ), 
        .C(\A_DOUT_TEMPR101[21] ), .D(\A_DOUT_TEMPR102[21] ), .Y(
        OR4_1700_Y));
    OR4 OR4_397 (.A(\A_DOUT_TEMPR12[27] ), .B(\A_DOUT_TEMPR13[27] ), 
        .C(\A_DOUT_TEMPR14[27] ), .D(\A_DOUT_TEMPR15[27] ), .Y(
        OR4_397_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%46%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R46C5 (
        .A_DOUT({nc21960, nc21961, nc21962, nc21963, nc21964, nc21965, 
        nc21966, nc21967, nc21968, nc21969, nc21970, nc21971, nc21972, 
        nc21973, nc21974, \A_DOUT_TEMPR46[29] , \A_DOUT_TEMPR46[28] , 
        \A_DOUT_TEMPR46[27] , \A_DOUT_TEMPR46[26] , 
        \A_DOUT_TEMPR46[25] }), .B_DOUT({nc21975, nc21976, nc21977, 
        nc21978, nc21979, nc21980, nc21981, nc21982, nc21983, nc21984, 
        nc21985, nc21986, nc21987, nc21988, nc21989, 
        \B_DOUT_TEMPR46[29] , \B_DOUT_TEMPR46[28] , 
        \B_DOUT_TEMPR46[27] , \B_DOUT_TEMPR46[26] , 
        \B_DOUT_TEMPR46[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[46][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%49%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R49C5 (
        .A_DOUT({nc21990, nc21991, nc21992, nc21993, nc21994, nc21995, 
        nc21996, nc21997, nc21998, nc21999, nc22000, nc22001, nc22002, 
        nc22003, nc22004, \A_DOUT_TEMPR49[29] , \A_DOUT_TEMPR49[28] , 
        \A_DOUT_TEMPR49[27] , \A_DOUT_TEMPR49[26] , 
        \A_DOUT_TEMPR49[25] }), .B_DOUT({nc22005, nc22006, nc22007, 
        nc22008, nc22009, nc22010, nc22011, nc22012, nc22013, nc22014, 
        nc22015, nc22016, nc22017, nc22018, nc22019, 
        \B_DOUT_TEMPR49[29] , \B_DOUT_TEMPR49[28] , 
        \B_DOUT_TEMPR49[27] , \B_DOUT_TEMPR49[26] , 
        \B_DOUT_TEMPR49[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%100%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R100C1 (
        .A_DOUT({nc22020, nc22021, nc22022, nc22023, nc22024, nc22025, 
        nc22026, nc22027, nc22028, nc22029, nc22030, nc22031, nc22032, 
        nc22033, nc22034, \A_DOUT_TEMPR100[9] , \A_DOUT_TEMPR100[8] , 
        \A_DOUT_TEMPR100[7] , \A_DOUT_TEMPR100[6] , 
        \A_DOUT_TEMPR100[5] }), .B_DOUT({nc22035, nc22036, nc22037, 
        nc22038, nc22039, nc22040, nc22041, nc22042, nc22043, nc22044, 
        nc22045, nc22046, nc22047, nc22048, nc22049, 
        \B_DOUT_TEMPR100[9] , \B_DOUT_TEMPR100[8] , 
        \B_DOUT_TEMPR100[7] , \B_DOUT_TEMPR100[6] , 
        \B_DOUT_TEMPR100[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[100][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1162 (.A(OR4_2774_Y), .B(OR4_2831_Y), .C(OR4_2365_Y), .D(
        OR4_1040_Y), .Y(OR4_1162_Y));
    OR4 OR4_2334 (.A(\A_DOUT_TEMPR75[4] ), .B(\A_DOUT_TEMPR76[4] ), .C(
        \A_DOUT_TEMPR77[4] ), .D(\A_DOUT_TEMPR78[4] ), .Y(OR4_2334_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%7%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R7C6 (
        .A_DOUT({nc22050, nc22051, nc22052, nc22053, nc22054, nc22055, 
        nc22056, nc22057, nc22058, nc22059, nc22060, nc22061, nc22062, 
        nc22063, nc22064, \A_DOUT_TEMPR7[34] , \A_DOUT_TEMPR7[33] , 
        \A_DOUT_TEMPR7[32] , \A_DOUT_TEMPR7[31] , \A_DOUT_TEMPR7[30] })
        , .B_DOUT({nc22065, nc22066, nc22067, nc22068, nc22069, 
        nc22070, nc22071, nc22072, nc22073, nc22074, nc22075, nc22076, 
        nc22077, nc22078, nc22079, \B_DOUT_TEMPR7[34] , 
        \B_DOUT_TEMPR7[33] , \B_DOUT_TEMPR7[32] , \B_DOUT_TEMPR7[31] , 
        \B_DOUT_TEMPR7[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_898 (.A(\B_DOUT_TEMPR4[29] ), .B(\B_DOUT_TEMPR5[29] ), .C(
        \B_DOUT_TEMPR6[29] ), .D(\B_DOUT_TEMPR7[29] ), .Y(OR4_898_Y));
    OR4 OR4_1711 (.A(\B_DOUT_TEMPR4[16] ), .B(\B_DOUT_TEMPR5[16] ), .C(
        \B_DOUT_TEMPR6[16] ), .D(\B_DOUT_TEMPR7[16] ), .Y(OR4_1711_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%51%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R51C6 (
        .A_DOUT({nc22080, nc22081, nc22082, nc22083, nc22084, nc22085, 
        nc22086, nc22087, nc22088, nc22089, nc22090, nc22091, nc22092, 
        nc22093, nc22094, \A_DOUT_TEMPR51[34] , \A_DOUT_TEMPR51[33] , 
        \A_DOUT_TEMPR51[32] , \A_DOUT_TEMPR51[31] , 
        \A_DOUT_TEMPR51[30] }), .B_DOUT({nc22095, nc22096, nc22097, 
        nc22098, nc22099, nc22100, nc22101, nc22102, nc22103, nc22104, 
        nc22105, nc22106, nc22107, nc22108, nc22109, 
        \B_DOUT_TEMPR51[34] , \B_DOUT_TEMPR51[33] , 
        \B_DOUT_TEMPR51[32] , \B_DOUT_TEMPR51[31] , 
        \B_DOUT_TEMPR51[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[51][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_691 (.A(\A_DOUT_TEMPR32[9] ), .B(\A_DOUT_TEMPR33[9] ), .C(
        \A_DOUT_TEMPR34[9] ), .D(\A_DOUT_TEMPR35[9] ), .Y(OR4_691_Y));
    OR4 OR4_854 (.A(\A_DOUT_TEMPR87[31] ), .B(\A_DOUT_TEMPR88[31] ), 
        .C(\A_DOUT_TEMPR89[31] ), .D(\A_DOUT_TEMPR90[31] ), .Y(
        OR4_854_Y));
    OR4 OR4_1334 (.A(\A_DOUT_TEMPR83[32] ), .B(\A_DOUT_TEMPR84[32] ), 
        .C(\A_DOUT_TEMPR85[32] ), .D(\A_DOUT_TEMPR86[32] ), .Y(
        OR4_1334_Y));
    OR4 OR4_552 (.A(\B_DOUT_TEMPR12[18] ), .B(\B_DOUT_TEMPR13[18] ), 
        .C(\B_DOUT_TEMPR14[18] ), .D(\B_DOUT_TEMPR15[18] ), .Y(
        OR4_552_Y));
    OR4 OR4_1658 (.A(\B_DOUT_TEMPR40[17] ), .B(\B_DOUT_TEMPR41[17] ), 
        .C(\B_DOUT_TEMPR42[17] ), .D(\B_DOUT_TEMPR43[17] ), .Y(
        OR4_1658_Y));
    OR4 OR4_49 (.A(OR4_449_Y), .B(OR4_1630_Y), .C(OR2_69_Y), .D(
        \B_DOUT_TEMPR74[13] ), .Y(OR4_49_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%92%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R92C2 (
        .A_DOUT({nc22110, nc22111, nc22112, nc22113, nc22114, nc22115, 
        nc22116, nc22117, nc22118, nc22119, nc22120, nc22121, nc22122, 
        nc22123, nc22124, \A_DOUT_TEMPR92[14] , \A_DOUT_TEMPR92[13] , 
        \A_DOUT_TEMPR92[12] , \A_DOUT_TEMPR92[11] , 
        \A_DOUT_TEMPR92[10] }), .B_DOUT({nc22125, nc22126, nc22127, 
        nc22128, nc22129, nc22130, nc22131, nc22132, nc22133, nc22134, 
        nc22135, nc22136, nc22137, nc22138, nc22139, 
        \B_DOUT_TEMPR92[14] , \B_DOUT_TEMPR92[13] , 
        \B_DOUT_TEMPR92[12] , \B_DOUT_TEMPR92[11] , 
        \B_DOUT_TEMPR92[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[92][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%6%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R6C7 (
        .A_DOUT({nc22140, nc22141, nc22142, nc22143, nc22144, nc22145, 
        nc22146, nc22147, nc22148, nc22149, nc22150, nc22151, nc22152, 
        nc22153, nc22154, \A_DOUT_TEMPR6[39] , \A_DOUT_TEMPR6[38] , 
        \A_DOUT_TEMPR6[37] , \A_DOUT_TEMPR6[36] , \A_DOUT_TEMPR6[35] })
        , .B_DOUT({nc22155, nc22156, nc22157, nc22158, nc22159, 
        nc22160, nc22161, nc22162, nc22163, nc22164, nc22165, nc22166, 
        nc22167, nc22168, nc22169, \B_DOUT_TEMPR6[39] , 
        \B_DOUT_TEMPR6[38] , \B_DOUT_TEMPR6[37] , \B_DOUT_TEMPR6[36] , 
        \B_DOUT_TEMPR6[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1870 (.A(\B_DOUT_TEMPR99[29] ), .B(\B_DOUT_TEMPR100[29] ), 
        .C(\B_DOUT_TEMPR101[29] ), .D(\B_DOUT_TEMPR102[29] ), .Y(
        OR4_1870_Y));
    OR4 OR4_494 (.A(OR4_541_Y), .B(OR4_343_Y), .C(OR2_6_Y), .D(
        \A_DOUT_TEMPR74[34] ), .Y(OR4_494_Y));
    OR4 OR4_2412 (.A(\A_DOUT_TEMPR83[21] ), .B(\A_DOUT_TEMPR84[21] ), 
        .C(\A_DOUT_TEMPR85[21] ), .D(\A_DOUT_TEMPR86[21] ), .Y(
        OR4_2412_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%112%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R112C5 (
        .A_DOUT({nc22170, nc22171, nc22172, nc22173, nc22174, nc22175, 
        nc22176, nc22177, nc22178, nc22179, nc22180, nc22181, nc22182, 
        nc22183, nc22184, \A_DOUT_TEMPR112[29] , \A_DOUT_TEMPR112[28] , 
        \A_DOUT_TEMPR112[27] , \A_DOUT_TEMPR112[26] , 
        \A_DOUT_TEMPR112[25] }), .B_DOUT({nc22185, nc22186, nc22187, 
        nc22188, nc22189, nc22190, nc22191, nc22192, nc22193, nc22194, 
        nc22195, nc22196, nc22197, nc22198, nc22199, 
        \B_DOUT_TEMPR112[29] , \B_DOUT_TEMPR112[28] , 
        \B_DOUT_TEMPR112[27] , \B_DOUT_TEMPR112[26] , 
        \B_DOUT_TEMPR112[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[112][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1307 (.A(OR4_2856_Y), .B(OR4_1451_Y), .C(OR4_842_Y), .D(
        OR4_147_Y), .Y(OR4_1307_Y));
    OR4 OR4_1202 (.A(OR4_1404_Y), .B(OR4_3026_Y), .C(OR4_606_Y), .D(
        OR4_2855_Y), .Y(OR4_1202_Y));
    OR4 OR4_2418 (.A(OR4_103_Y), .B(OR4_1049_Y), .C(OR4_676_Y), .D(
        OR4_2151_Y), .Y(OR4_2418_Y));
    OR4 OR4_1874 (.A(OR4_2555_Y), .B(OR4_2359_Y), .C(OR2_54_Y), .D(
        \B_DOUT_TEMPR74[38] ), .Y(OR4_1874_Y));
    OR4 OR4_2751 (.A(\B_DOUT_TEMPR36[24] ), .B(\B_DOUT_TEMPR37[24] ), 
        .C(\B_DOUT_TEMPR38[24] ), .D(\B_DOUT_TEMPR39[24] ), .Y(
        OR4_2751_Y));
    OR4 OR4_338 (.A(\B_DOUT_TEMPR4[20] ), .B(\B_DOUT_TEMPR5[20] ), .C(
        \B_DOUT_TEMPR6[20] ), .D(\B_DOUT_TEMPR7[20] ), .Y(OR4_338_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%0%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R0C7 (
        .A_DOUT({nc22200, nc22201, nc22202, nc22203, nc22204, nc22205, 
        nc22206, nc22207, nc22208, nc22209, nc22210, nc22211, nc22212, 
        nc22213, nc22214, \A_DOUT_TEMPR0[39] , \A_DOUT_TEMPR0[38] , 
        \A_DOUT_TEMPR0[37] , \A_DOUT_TEMPR0[36] , \A_DOUT_TEMPR0[35] })
        , .B_DOUT({nc22215, nc22216, nc22217, nc22218, nc22219, 
        nc22220, nc22221, nc22222, nc22223, nc22224, nc22225, nc22226, 
        nc22227, nc22228, nc22229, \B_DOUT_TEMPR0[39] , 
        \B_DOUT_TEMPR0[38] , \B_DOUT_TEMPR0[37] , \B_DOUT_TEMPR0[36] , 
        \B_DOUT_TEMPR0[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1188 (.A(\B_DOUT_TEMPR16[37] ), .B(\B_DOUT_TEMPR17[37] ), 
        .C(\B_DOUT_TEMPR18[37] ), .D(\B_DOUT_TEMPR19[37] ), .Y(
        OR4_1188_Y));
    OR4 OR4_1898 (.A(\A_DOUT_TEMPR44[2] ), .B(\A_DOUT_TEMPR45[2] ), .C(
        \A_DOUT_TEMPR46[2] ), .D(\A_DOUT_TEMPR47[2] ), .Y(OR4_1898_Y));
    OR4 OR4_1020 (.A(\A_DOUT_TEMPR8[0] ), .B(\A_DOUT_TEMPR9[0] ), .C(
        \A_DOUT_TEMPR10[0] ), .D(\A_DOUT_TEMPR11[0] ), .Y(OR4_1020_Y));
    OR4 OR4_735 (.A(\A_DOUT_TEMPR75[3] ), .B(\A_DOUT_TEMPR76[3] ), .C(
        \A_DOUT_TEMPR77[3] ), .D(\A_DOUT_TEMPR78[3] ), .Y(OR4_735_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%58%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R58C2 (
        .A_DOUT({nc22230, nc22231, nc22232, nc22233, nc22234, nc22235, 
        nc22236, nc22237, nc22238, nc22239, nc22240, nc22241, nc22242, 
        nc22243, nc22244, \A_DOUT_TEMPR58[14] , \A_DOUT_TEMPR58[13] , 
        \A_DOUT_TEMPR58[12] , \A_DOUT_TEMPR58[11] , 
        \A_DOUT_TEMPR58[10] }), .B_DOUT({nc22245, nc22246, nc22247, 
        nc22248, nc22249, nc22250, nc22251, nc22252, nc22253, nc22254, 
        nc22255, nc22256, nc22257, nc22258, nc22259, 
        \B_DOUT_TEMPR58[14] , \B_DOUT_TEMPR58[13] , 
        \B_DOUT_TEMPR58[12] , \B_DOUT_TEMPR58[11] , 
        \B_DOUT_TEMPR58[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[58][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%93%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R93C1 (
        .A_DOUT({nc22260, nc22261, nc22262, nc22263, nc22264, nc22265, 
        nc22266, nc22267, nc22268, nc22269, nc22270, nc22271, nc22272, 
        nc22273, nc22274, \A_DOUT_TEMPR93[9] , \A_DOUT_TEMPR93[8] , 
        \A_DOUT_TEMPR93[7] , \A_DOUT_TEMPR93[6] , \A_DOUT_TEMPR93[5] })
        , .B_DOUT({nc22275, nc22276, nc22277, nc22278, nc22279, 
        nc22280, nc22281, nc22282, nc22283, nc22284, nc22285, nc22286, 
        nc22287, nc22288, nc22289, \B_DOUT_TEMPR93[9] , 
        \B_DOUT_TEMPR93[8] , \B_DOUT_TEMPR93[7] , \B_DOUT_TEMPR93[6] , 
        \B_DOUT_TEMPR93[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[93][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1413 (.A(\B_DOUT_TEMPR36[34] ), .B(\B_DOUT_TEMPR37[34] ), 
        .C(\B_DOUT_TEMPR38[34] ), .D(\B_DOUT_TEMPR39[34] ), .Y(
        OR4_1413_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%32%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R32C0 (
        .A_DOUT({nc22290, nc22291, nc22292, nc22293, nc22294, nc22295, 
        nc22296, nc22297, nc22298, nc22299, nc22300, nc22301, nc22302, 
        nc22303, nc22304, \A_DOUT_TEMPR32[4] , \A_DOUT_TEMPR32[3] , 
        \A_DOUT_TEMPR32[2] , \A_DOUT_TEMPR32[1] , \A_DOUT_TEMPR32[0] })
        , .B_DOUT({nc22305, nc22306, nc22307, nc22308, nc22309, 
        nc22310, nc22311, nc22312, nc22313, nc22314, nc22315, nc22316, 
        nc22317, nc22318, nc22319, \B_DOUT_TEMPR32[4] , 
        \B_DOUT_TEMPR32[3] , \B_DOUT_TEMPR32[2] , \B_DOUT_TEMPR32[1] , 
        \B_DOUT_TEMPR32[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[32][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%28%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R28C1 (
        .A_DOUT({nc22320, nc22321, nc22322, nc22323, nc22324, nc22325, 
        nc22326, nc22327, nc22328, nc22329, nc22330, nc22331, nc22332, 
        nc22333, nc22334, \A_DOUT_TEMPR28[9] , \A_DOUT_TEMPR28[8] , 
        \A_DOUT_TEMPR28[7] , \A_DOUT_TEMPR28[6] , \A_DOUT_TEMPR28[5] })
        , .B_DOUT({nc22335, nc22336, nc22337, nc22338, nc22339, 
        nc22340, nc22341, nc22342, nc22343, nc22344, nc22345, nc22346, 
        nc22347, nc22348, nc22349, \B_DOUT_TEMPR28[9] , 
        \B_DOUT_TEMPR28[8] , \B_DOUT_TEMPR28[7] , \B_DOUT_TEMPR28[6] , 
        \B_DOUT_TEMPR28[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    CFG3 #( .INIT(8'h80) )  CFG3_9 (.A(B_BLK_EN), .B(B_ADDR[18]), .C(
        B_ADDR[17]), .Y(CFG3_9_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%87%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R87C4 (
        .A_DOUT({nc22350, nc22351, nc22352, nc22353, nc22354, nc22355, 
        nc22356, nc22357, nc22358, nc22359, nc22360, nc22361, nc22362, 
        nc22363, nc22364, \A_DOUT_TEMPR87[24] , \A_DOUT_TEMPR87[23] , 
        \A_DOUT_TEMPR87[22] , \A_DOUT_TEMPR87[21] , 
        \A_DOUT_TEMPR87[20] }), .B_DOUT({nc22365, nc22366, nc22367, 
        nc22368, nc22369, nc22370, nc22371, nc22372, nc22373, nc22374, 
        nc22375, nc22376, nc22377, nc22378, nc22379, 
        \B_DOUT_TEMPR87[24] , \B_DOUT_TEMPR87[23] , 
        \B_DOUT_TEMPR87[22] , \B_DOUT_TEMPR87[21] , 
        \B_DOUT_TEMPR87[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[87][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_11 (.A(OR4_2944_Y), .B(OR4_705_Y), .C(OR2_72_Y), .D(
        \A_DOUT_TEMPR74[26] ), .Y(OR4_11_Y));
    OR4 OR4_719 (.A(\B_DOUT_TEMPR56[23] ), .B(\B_DOUT_TEMPR57[23] ), 
        .C(\B_DOUT_TEMPR58[23] ), .D(\B_DOUT_TEMPR59[23] ), .Y(
        OR4_719_Y));
    OR4 OR4_58 (.A(OR4_1720_Y), .B(OR4_2548_Y), .C(OR4_1605_Y), .D(
        OR4_2366_Y), .Y(OR4_58_Y));
    OR4 OR4_2941 (.A(\A_DOUT_TEMPR0[0] ), .B(\A_DOUT_TEMPR1[0] ), .C(
        \A_DOUT_TEMPR2[0] ), .D(\A_DOUT_TEMPR3[0] ), .Y(OR4_2941_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%28%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R28C7 (
        .A_DOUT({nc22380, nc22381, nc22382, nc22383, nc22384, nc22385, 
        nc22386, nc22387, nc22388, nc22389, nc22390, nc22391, nc22392, 
        nc22393, nc22394, \A_DOUT_TEMPR28[39] , \A_DOUT_TEMPR28[38] , 
        \A_DOUT_TEMPR28[37] , \A_DOUT_TEMPR28[36] , 
        \A_DOUT_TEMPR28[35] }), .B_DOUT({nc22395, nc22396, nc22397, 
        nc22398, nc22399, nc22400, nc22401, nc22402, nc22403, nc22404, 
        nc22405, nc22406, nc22407, nc22408, nc22409, 
        \B_DOUT_TEMPR28[39] , \B_DOUT_TEMPR28[38] , 
        \B_DOUT_TEMPR28[37] , \B_DOUT_TEMPR28[36] , 
        \B_DOUT_TEMPR28[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2510 (.A(OR4_2043_Y), .B(OR4_2878_Y), .C(OR2_46_Y), .D(
        \B_DOUT_TEMPR74[25] ), .Y(OR4_2510_Y));
    OR4 OR4_1404 (.A(\B_DOUT_TEMPR32[21] ), .B(\B_DOUT_TEMPR33[21] ), 
        .C(\B_DOUT_TEMPR34[21] ), .D(\B_DOUT_TEMPR35[21] ), .Y(
        OR4_1404_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%79%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R79C3 (
        .A_DOUT({nc22410, nc22411, nc22412, nc22413, nc22414, nc22415, 
        nc22416, nc22417, nc22418, nc22419, nc22420, nc22421, nc22422, 
        nc22423, nc22424, \A_DOUT_TEMPR79[19] , \A_DOUT_TEMPR79[18] , 
        \A_DOUT_TEMPR79[17] , \A_DOUT_TEMPR79[16] , 
        \A_DOUT_TEMPR79[15] }), .B_DOUT({nc22425, nc22426, nc22427, 
        nc22428, nc22429, nc22430, nc22431, nc22432, nc22433, nc22434, 
        nc22435, nc22436, nc22437, nc22438, nc22439, 
        \B_DOUT_TEMPR79[19] , \B_DOUT_TEMPR79[18] , 
        \B_DOUT_TEMPR79[17] , \B_DOUT_TEMPR79[16] , 
        \B_DOUT_TEMPR79[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[79][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[20]  (.A(OR4_1761_Y), .B(OR4_1220_Y), .C(OR4_935_Y)
        , .D(OR4_2401_Y), .Y(B_DOUT[20]));
    OR4 OR4_2395 (.A(OR4_1169_Y), .B(OR4_2327_Y), .C(OR2_11_Y), .D(
        \A_DOUT_TEMPR74[14] ), .Y(OR4_2395_Y));
    OR4 OR4_1883 (.A(\B_DOUT_TEMPR16[19] ), .B(\B_DOUT_TEMPR17[19] ), 
        .C(\B_DOUT_TEMPR18[19] ), .D(\B_DOUT_TEMPR19[19] ), .Y(
        OR4_1883_Y));
    OR4 OR4_615 (.A(\A_DOUT_TEMPR16[30] ), .B(\A_DOUT_TEMPR17[30] ), 
        .C(\A_DOUT_TEMPR18[30] ), .D(\A_DOUT_TEMPR19[30] ), .Y(
        OR4_615_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%13%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R13C3 (
        .A_DOUT({nc22440, nc22441, nc22442, nc22443, nc22444, nc22445, 
        nc22446, nc22447, nc22448, nc22449, nc22450, nc22451, nc22452, 
        nc22453, nc22454, \A_DOUT_TEMPR13[19] , \A_DOUT_TEMPR13[18] , 
        \A_DOUT_TEMPR13[17] , \A_DOUT_TEMPR13[16] , 
        \A_DOUT_TEMPR13[15] }), .B_DOUT({nc22455, nc22456, nc22457, 
        nc22458, nc22459, nc22460, nc22461, nc22462, nc22463, nc22464, 
        nc22465, nc22466, nc22467, nc22468, nc22469, 
        \B_DOUT_TEMPR13[19] , \B_DOUT_TEMPR13[18] , 
        \B_DOUT_TEMPR13[17] , \B_DOUT_TEMPR13[16] , 
        \B_DOUT_TEMPR13[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%31%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R31C6 (
        .A_DOUT({nc22470, nc22471, nc22472, nc22473, nc22474, nc22475, 
        nc22476, nc22477, nc22478, nc22479, nc22480, nc22481, nc22482, 
        nc22483, nc22484, \A_DOUT_TEMPR31[34] , \A_DOUT_TEMPR31[33] , 
        \A_DOUT_TEMPR31[32] , \A_DOUT_TEMPR31[31] , 
        \A_DOUT_TEMPR31[30] }), .B_DOUT({nc22485, nc22486, nc22487, 
        nc22488, nc22489, nc22490, nc22491, nc22492, nc22493, nc22494, 
        nc22495, nc22496, nc22497, nc22498, nc22499, 
        \B_DOUT_TEMPR31[34] , \B_DOUT_TEMPR31[33] , 
        \B_DOUT_TEMPR31[32] , \B_DOUT_TEMPR31[31] , 
        \B_DOUT_TEMPR31[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_427 (.A(\A_DOUT_TEMPR107[8] ), .B(\A_DOUT_TEMPR108[8] ), 
        .C(\A_DOUT_TEMPR109[8] ), .D(\A_DOUT_TEMPR110[8] ), .Y(
        OR4_427_Y));
    OR4 OR4_2967 (.A(\B_DOUT_TEMPR0[30] ), .B(\B_DOUT_TEMPR1[30] ), .C(
        \B_DOUT_TEMPR2[30] ), .D(\B_DOUT_TEMPR3[30] ), .Y(OR4_2967_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%15%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R15C3 (
        .A_DOUT({nc22500, nc22501, nc22502, nc22503, nc22504, nc22505, 
        nc22506, nc22507, nc22508, nc22509, nc22510, nc22511, nc22512, 
        nc22513, nc22514, \A_DOUT_TEMPR15[19] , \A_DOUT_TEMPR15[18] , 
        \A_DOUT_TEMPR15[17] , \A_DOUT_TEMPR15[16] , 
        \A_DOUT_TEMPR15[15] }), .B_DOUT({nc22515, nc22516, nc22517, 
        nc22518, nc22519, nc22520, nc22521, nc22522, nc22523, nc22524, 
        nc22525, nc22526, nc22527, nc22528, nc22529, 
        \B_DOUT_TEMPR15[19] , \B_DOUT_TEMPR15[18] , 
        \B_DOUT_TEMPR15[17] , \B_DOUT_TEMPR15[16] , 
        \B_DOUT_TEMPR15[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[15][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_219 (.A(OR4_2116_Y), .B(OR4_1931_Y), .C(OR4_2815_Y), .D(
        OR4_972_Y), .Y(OR4_219_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%58%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R58C3 (
        .A_DOUT({nc22530, nc22531, nc22532, nc22533, nc22534, nc22535, 
        nc22536, nc22537, nc22538, nc22539, nc22540, nc22541, nc22542, 
        nc22543, nc22544, \A_DOUT_TEMPR58[19] , \A_DOUT_TEMPR58[18] , 
        \A_DOUT_TEMPR58[17] , \A_DOUT_TEMPR58[16] , 
        \A_DOUT_TEMPR58[15] }), .B_DOUT({nc22545, nc22546, nc22547, 
        nc22548, nc22549, nc22550, nc22551, nc22552, nc22553, nc22554, 
        nc22555, nc22556, nc22557, nc22558, nc22559, 
        \B_DOUT_TEMPR58[19] , \B_DOUT_TEMPR58[18] , 
        \B_DOUT_TEMPR58[17] , \B_DOUT_TEMPR58[16] , 
        \B_DOUT_TEMPR58[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[58][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_938 (.A(\A_DOUT_TEMPR4[19] ), .B(\A_DOUT_TEMPR5[19] ), .C(
        \A_DOUT_TEMPR6[19] ), .D(\A_DOUT_TEMPR7[19] ), .Y(OR4_938_Y));
    OR4 OR4_1789 (.A(\A_DOUT_TEMPR79[11] ), .B(\A_DOUT_TEMPR80[11] ), 
        .C(\A_DOUT_TEMPR81[11] ), .D(\A_DOUT_TEMPR82[11] ), .Y(
        OR4_1789_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%83%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R83C6 (
        .A_DOUT({nc22560, nc22561, nc22562, nc22563, nc22564, nc22565, 
        nc22566, nc22567, nc22568, nc22569, nc22570, nc22571, nc22572, 
        nc22573, nc22574, \A_DOUT_TEMPR83[34] , \A_DOUT_TEMPR83[33] , 
        \A_DOUT_TEMPR83[32] , \A_DOUT_TEMPR83[31] , 
        \A_DOUT_TEMPR83[30] }), .B_DOUT({nc22575, nc22576, nc22577, 
        nc22578, nc22579, nc22580, nc22581, nc22582, nc22583, nc22584, 
        nc22585, nc22586, nc22587, nc22588, nc22589, 
        \B_DOUT_TEMPR83[34] , \B_DOUT_TEMPR83[33] , 
        \B_DOUT_TEMPR83[32] , \B_DOUT_TEMPR83[31] , 
        \B_DOUT_TEMPR83[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[83][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2430 (.A(\B_DOUT_TEMPR79[28] ), .B(\B_DOUT_TEMPR80[28] ), 
        .C(\B_DOUT_TEMPR81[28] ), .D(\B_DOUT_TEMPR82[28] ), .Y(
        OR4_2430_Y));
    OR4 OR4_2453 (.A(\A_DOUT_TEMPR0[25] ), .B(\A_DOUT_TEMPR1[25] ), .C(
        \A_DOUT_TEMPR2[25] ), .D(\A_DOUT_TEMPR3[25] ), .Y(OR4_2453_Y));
    OR4 OR4_713 (.A(\A_DOUT_TEMPR56[20] ), .B(\A_DOUT_TEMPR57[20] ), 
        .C(\A_DOUT_TEMPR58[20] ), .D(\A_DOUT_TEMPR59[20] ), .Y(
        OR4_713_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%54%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R54C1 (
        .A_DOUT({nc22590, nc22591, nc22592, nc22593, nc22594, nc22595, 
        nc22596, nc22597, nc22598, nc22599, nc22600, nc22601, nc22602, 
        nc22603, nc22604, \A_DOUT_TEMPR54[9] , \A_DOUT_TEMPR54[8] , 
        \A_DOUT_TEMPR54[7] , \A_DOUT_TEMPR54[6] , \A_DOUT_TEMPR54[5] })
        , .B_DOUT({nc22605, nc22606, nc22607, nc22608, nc22609, 
        nc22610, nc22611, nc22612, nc22613, nc22614, nc22615, nc22616, 
        nc22617, nc22618, nc22619, \B_DOUT_TEMPR54[9] , 
        \B_DOUT_TEMPR54[8] , \B_DOUT_TEMPR54[7] , \B_DOUT_TEMPR54[6] , 
        \B_DOUT_TEMPR54[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[54][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1430 (.A(OR4_252_Y), .B(OR4_1444_Y), .C(OR4_2494_Y), .D(
        OR4_697_Y), .Y(OR4_1430_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%50%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R50C4 (
        .A_DOUT({nc22620, nc22621, nc22622, nc22623, nc22624, nc22625, 
        nc22626, nc22627, nc22628, nc22629, nc22630, nc22631, nc22632, 
        nc22633, nc22634, \A_DOUT_TEMPR50[24] , \A_DOUT_TEMPR50[23] , 
        \A_DOUT_TEMPR50[22] , \A_DOUT_TEMPR50[21] , 
        \A_DOUT_TEMPR50[20] }), .B_DOUT({nc22635, nc22636, nc22637, 
        nc22638, nc22639, nc22640, nc22641, nc22642, nc22643, nc22644, 
        nc22645, nc22646, nc22647, nc22648, nc22649, 
        \B_DOUT_TEMPR50[24] , \B_DOUT_TEMPR50[23] , 
        \B_DOUT_TEMPR50[22] , \B_DOUT_TEMPR50[21] , 
        \B_DOUT_TEMPR50[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2128 (.A(\B_DOUT_TEMPR79[39] ), .B(\B_DOUT_TEMPR80[39] ), 
        .C(\B_DOUT_TEMPR81[39] ), .D(\B_DOUT_TEMPR82[39] ), .Y(
        OR4_2128_Y));
    OR4 OR4_2879 (.A(OR4_438_Y), .B(OR4_247_Y), .C(OR4_192_Y), .D(
        OR4_892_Y), .Y(OR4_2879_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%77%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R77C3 (
        .A_DOUT({nc22650, nc22651, nc22652, nc22653, nc22654, nc22655, 
        nc22656, nc22657, nc22658, nc22659, nc22660, nc22661, nc22662, 
        nc22663, nc22664, \A_DOUT_TEMPR77[19] , \A_DOUT_TEMPR77[18] , 
        \A_DOUT_TEMPR77[17] , \A_DOUT_TEMPR77[16] , 
        \A_DOUT_TEMPR77[15] }), .B_DOUT({nc22665, nc22666, nc22667, 
        nc22668, nc22669, nc22670, nc22671, nc22672, nc22673, nc22674, 
        nc22675, nc22676, nc22677, nc22678, nc22679, 
        \B_DOUT_TEMPR77[19] , \B_DOUT_TEMPR77[18] , 
        \B_DOUT_TEMPR77[17] , \B_DOUT_TEMPR77[16] , 
        \B_DOUT_TEMPR77[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[77][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%0%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R0C0 (
        .A_DOUT({nc22680, nc22681, nc22682, nc22683, nc22684, nc22685, 
        nc22686, nc22687, nc22688, nc22689, nc22690, nc22691, nc22692, 
        nc22693, nc22694, \A_DOUT_TEMPR0[4] , \A_DOUT_TEMPR0[3] , 
        \A_DOUT_TEMPR0[2] , \A_DOUT_TEMPR0[1] , \A_DOUT_TEMPR0[0] }), 
        .B_DOUT({nc22695, nc22696, nc22697, nc22698, nc22699, nc22700, 
        nc22701, nc22702, nc22703, nc22704, nc22705, nc22706, nc22707, 
        nc22708, nc22709, \B_DOUT_TEMPR0[4] , \B_DOUT_TEMPR0[3] , 
        \B_DOUT_TEMPR0[2] , \B_DOUT_TEMPR0[1] , \B_DOUT_TEMPR0[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[0][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[0] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%60%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R60C7 (
        .A_DOUT({nc22710, nc22711, nc22712, nc22713, nc22714, nc22715, 
        nc22716, nc22717, nc22718, nc22719, nc22720, nc22721, nc22722, 
        nc22723, nc22724, \A_DOUT_TEMPR60[39] , \A_DOUT_TEMPR60[38] , 
        \A_DOUT_TEMPR60[37] , \A_DOUT_TEMPR60[36] , 
        \A_DOUT_TEMPR60[35] }), .B_DOUT({nc22725, nc22726, nc22727, 
        nc22728, nc22729, nc22730, nc22731, nc22732, nc22733, nc22734, 
        nc22735, nc22736, nc22737, nc22738, nc22739, 
        \B_DOUT_TEMPR60[39] , \B_DOUT_TEMPR60[38] , 
        \B_DOUT_TEMPR60[37] , \B_DOUT_TEMPR60[36] , 
        \B_DOUT_TEMPR60[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[60][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1186 (.A(OR4_2705_Y), .B(OR4_1698_Y), .C(OR4_1917_Y), .D(
        OR4_1708_Y), .Y(OR4_1186_Y));
    OR4 OR4_2385 (.A(\A_DOUT_TEMPR95[3] ), .B(\A_DOUT_TEMPR96[3] ), .C(
        \A_DOUT_TEMPR97[3] ), .D(\A_DOUT_TEMPR98[3] ), .Y(OR4_2385_Y));
    OR4 OR4_1426 (.A(\A_DOUT_TEMPR87[3] ), .B(\A_DOUT_TEMPR88[3] ), .C(
        \A_DOUT_TEMPR89[3] ), .D(\A_DOUT_TEMPR90[3] ), .Y(OR4_1426_Y));
    OR4 OR4_2243 (.A(OR4_2462_Y), .B(OR4_316_Y), .C(OR4_1047_Y), .D(
        OR4_1334_Y), .Y(OR4_2243_Y));
    OR4 OR4_1741 (.A(\A_DOUT_TEMPR99[6] ), .B(\A_DOUT_TEMPR100[6] ), 
        .C(\A_DOUT_TEMPR101[6] ), .D(\A_DOUT_TEMPR102[6] ), .Y(
        OR4_1741_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%107%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R107C7 (
        .A_DOUT({nc22740, nc22741, nc22742, nc22743, nc22744, nc22745, 
        nc22746, nc22747, nc22748, nc22749, nc22750, nc22751, nc22752, 
        nc22753, nc22754, \A_DOUT_TEMPR107[39] , \A_DOUT_TEMPR107[38] , 
        \A_DOUT_TEMPR107[37] , \A_DOUT_TEMPR107[36] , 
        \A_DOUT_TEMPR107[35] }), .B_DOUT({nc22755, nc22756, nc22757, 
        nc22758, nc22759, nc22760, nc22761, nc22762, nc22763, nc22764, 
        nc22765, nc22766, nc22767, nc22768, nc22769, 
        \B_DOUT_TEMPR107[39] , \B_DOUT_TEMPR107[38] , 
        \B_DOUT_TEMPR107[37] , \B_DOUT_TEMPR107[36] , 
        \B_DOUT_TEMPR107[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[107][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1269 (.A(\A_DOUT_TEMPR99[16] ), .B(\A_DOUT_TEMPR100[16] ), 
        .C(\A_DOUT_TEMPR101[16] ), .D(\A_DOUT_TEMPR102[16] ), .Y(
        OR4_1269_Y));
    OR4 OR4_1588 (.A(\B_DOUT_TEMPR16[24] ), .B(\B_DOUT_TEMPR17[24] ), 
        .C(\B_DOUT_TEMPR18[24] ), .D(\B_DOUT_TEMPR19[24] ), .Y(
        OR4_1588_Y));
    OR4 OR4_138 (.A(\A_DOUT_TEMPR28[24] ), .B(\A_DOUT_TEMPR29[24] ), 
        .C(\A_DOUT_TEMPR30[24] ), .D(\A_DOUT_TEMPR31[24] ), .Y(
        OR4_138_Y));
    OR4 OR4_2235 (.A(\A_DOUT_TEMPR91[12] ), .B(\A_DOUT_TEMPR92[12] ), 
        .C(\A_DOUT_TEMPR93[12] ), .D(\A_DOUT_TEMPR94[12] ), .Y(
        OR4_2235_Y));
    OR4 OR4_1798 (.A(\B_DOUT_TEMPR75[28] ), .B(\B_DOUT_TEMPR76[28] ), 
        .C(\B_DOUT_TEMPR77[28] ), .D(\B_DOUT_TEMPR78[28] ), .Y(
        OR4_1798_Y));
    OR4 OR4_2860 (.A(\A_DOUT_TEMPR32[31] ), .B(\A_DOUT_TEMPR33[31] ), 
        .C(\A_DOUT_TEMPR34[31] ), .D(\A_DOUT_TEMPR35[31] ), .Y(
        OR4_2860_Y));
    OR4 OR4_218 (.A(\B_DOUT_TEMPR0[5] ), .B(\B_DOUT_TEMPR1[5] ), .C(
        \B_DOUT_TEMPR2[5] ), .D(\B_DOUT_TEMPR3[5] ), .Y(OR4_218_Y));
    OR4 OR4_2308 (.A(OR4_656_Y), .B(OR4_973_Y), .C(OR4_2549_Y), .D(
        OR4_425_Y), .Y(OR4_2308_Y));
    OR2 OR2_58 (.A(\A_DOUT_TEMPR72[4] ), .B(\A_DOUT_TEMPR73[4] ), .Y(
        OR2_58_Y));
    OR4 OR4_339 (.A(\B_DOUT_TEMPR103[9] ), .B(\B_DOUT_TEMPR104[9] ), 
        .C(\B_DOUT_TEMPR105[9] ), .D(\B_DOUT_TEMPR106[9] ), .Y(
        OR4_339_Y));
    OR4 OR4_2171 (.A(\A_DOUT_TEMPR4[34] ), .B(\A_DOUT_TEMPR5[34] ), .C(
        \A_DOUT_TEMPR6[34] ), .D(\A_DOUT_TEMPR7[34] ), .Y(OR4_2171_Y));
    OR4 OR4_894 (.A(\B_DOUT_TEMPR111[6] ), .B(\B_DOUT_TEMPR112[6] ), 
        .C(\B_DOUT_TEMPR113[6] ), .D(\B_DOUT_TEMPR114[6] ), .Y(
        OR4_894_Y));
    OR4 OR4_2915 (.A(OR4_2528_Y), .B(OR4_2323_Y), .C(OR4_2267_Y), .D(
        OR4_1941_Y), .Y(OR4_2915_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%10%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R10C1 (
        .A_DOUT({nc22770, nc22771, nc22772, nc22773, nc22774, nc22775, 
        nc22776, nc22777, nc22778, nc22779, nc22780, nc22781, nc22782, 
        nc22783, nc22784, \A_DOUT_TEMPR10[9] , \A_DOUT_TEMPR10[8] , 
        \A_DOUT_TEMPR10[7] , \A_DOUT_TEMPR10[6] , \A_DOUT_TEMPR10[5] })
        , .B_DOUT({nc22785, nc22786, nc22787, nc22788, nc22789, 
        nc22790, nc22791, nc22792, nc22793, nc22794, nc22795, nc22796, 
        nc22797, nc22798, nc22799, \B_DOUT_TEMPR10[9] , 
        \B_DOUT_TEMPR10[8] , \B_DOUT_TEMPR10[7] , \B_DOUT_TEMPR10[6] , 
        \B_DOUT_TEMPR10[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1235 (.A(OR4_1101_Y), .B(OR4_1808_Y), .C(OR4_1021_Y), .D(
        OR4_2983_Y), .Y(OR4_1235_Y));
    OR4 OR4_2823 (.A(\A_DOUT_TEMPR12[11] ), .B(\A_DOUT_TEMPR13[11] ), 
        .C(\A_DOUT_TEMPR14[11] ), .D(\A_DOUT_TEMPR15[11] ), .Y(
        OR4_2823_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%38%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R38C2 (
        .A_DOUT({nc22800, nc22801, nc22802, nc22803, nc22804, nc22805, 
        nc22806, nc22807, nc22808, nc22809, nc22810, nc22811, nc22812, 
        nc22813, nc22814, \A_DOUT_TEMPR38[14] , \A_DOUT_TEMPR38[13] , 
        \A_DOUT_TEMPR38[12] , \A_DOUT_TEMPR38[11] , 
        \A_DOUT_TEMPR38[10] }), .B_DOUT({nc22815, nc22816, nc22817, 
        nc22818, nc22819, nc22820, nc22821, nc22822, nc22823, nc22824, 
        nc22825, nc22826, nc22827, nc22828, nc22829, 
        \B_DOUT_TEMPR38[14] , \B_DOUT_TEMPR38[13] , 
        \B_DOUT_TEMPR38[12] , \B_DOUT_TEMPR38[11] , 
        \B_DOUT_TEMPR38[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[38][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_592 (.A(\B_DOUT_TEMPR107[8] ), .B(\B_DOUT_TEMPR108[8] ), 
        .C(\B_DOUT_TEMPR109[8] ), .D(\B_DOUT_TEMPR110[8] ), .Y(
        OR4_592_Y));
    OR4 OR4_1859 (.A(\A_DOUT_TEMPR68[32] ), .B(\A_DOUT_TEMPR69[32] ), 
        .C(\A_DOUT_TEMPR70[32] ), .D(\A_DOUT_TEMPR71[32] ), .Y(
        OR4_1859_Y));
    OR4 OR4_2864 (.A(\B_DOUT_TEMPR107[13] ), .B(\B_DOUT_TEMPR108[13] ), 
        .C(\B_DOUT_TEMPR109[13] ), .D(\B_DOUT_TEMPR110[13] ), .Y(
        OR4_2864_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%21%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R21C1 (
        .A_DOUT({nc22830, nc22831, nc22832, nc22833, nc22834, nc22835, 
        nc22836, nc22837, nc22838, nc22839, nc22840, nc22841, nc22842, 
        nc22843, nc22844, \A_DOUT_TEMPR21[9] , \A_DOUT_TEMPR21[8] , 
        \A_DOUT_TEMPR21[7] , \A_DOUT_TEMPR21[6] , \A_DOUT_TEMPR21[5] })
        , .B_DOUT({nc22845, nc22846, nc22847, nc22848, nc22849, 
        nc22850, nc22851, nc22852, nc22853, nc22854, nc22855, nc22856, 
        nc22857, nc22858, nc22859, \B_DOUT_TEMPR21[9] , 
        \B_DOUT_TEMPR21[8] , \B_DOUT_TEMPR21[7] , \B_DOUT_TEMPR21[6] , 
        \B_DOUT_TEMPR21[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%4%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R4C0 (
        .A_DOUT({nc22860, nc22861, nc22862, nc22863, nc22864, nc22865, 
        nc22866, nc22867, nc22868, nc22869, nc22870, nc22871, nc22872, 
        nc22873, nc22874, \A_DOUT_TEMPR4[4] , \A_DOUT_TEMPR4[3] , 
        \A_DOUT_TEMPR4[2] , \A_DOUT_TEMPR4[1] , \A_DOUT_TEMPR4[0] }), 
        .B_DOUT({nc22875, nc22876, nc22877, nc22878, nc22879, nc22880, 
        nc22881, nc22882, nc22883, nc22884, nc22885, nc22886, nc22887, 
        nc22888, nc22889, \B_DOUT_TEMPR4[4] , \B_DOUT_TEMPR4[3] , 
        \B_DOUT_TEMPR4[2] , \B_DOUT_TEMPR4[1] , \B_DOUT_TEMPR4[0] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[4][0] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[1] , \BLKX1[0] , \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[4], A_DIN[3], A_DIN[2], A_DIN[1], 
        A_DIN[0]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[0] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], B_DIN[1], 
        B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1725 (.A(\B_DOUT_TEMPR32[5] ), .B(\B_DOUT_TEMPR33[5] ), .C(
        \B_DOUT_TEMPR34[5] ), .D(\B_DOUT_TEMPR35[5] ), .Y(OR4_1725_Y));
    OR4 OR4_2075 (.A(\A_DOUT_TEMPR40[34] ), .B(\A_DOUT_TEMPR41[34] ), 
        .C(\A_DOUT_TEMPR42[34] ), .D(\A_DOUT_TEMPR43[34] ), .Y(
        OR4_2075_Y));
    OR4 OR4_2619 (.A(\A_DOUT_TEMPR91[29] ), .B(\A_DOUT_TEMPR92[29] ), 
        .C(\A_DOUT_TEMPR93[29] ), .D(\A_DOUT_TEMPR94[29] ), .Y(
        OR4_2619_Y));
    OR4 OR4_2729 (.A(\A_DOUT_TEMPR75[15] ), .B(\A_DOUT_TEMPR76[15] ), 
        .C(\A_DOUT_TEMPR77[15] ), .D(\A_DOUT_TEMPR78[15] ), .Y(
        OR4_2729_Y));
    OR4 OR4_1204 (.A(\B_DOUT_TEMPR79[38] ), .B(\B_DOUT_TEMPR80[38] ), 
        .C(\B_DOUT_TEMPR81[38] ), .D(\B_DOUT_TEMPR82[38] ), .Y(
        OR4_1204_Y));
    OR4 OR4_1151 (.A(\B_DOUT_TEMPR99[1] ), .B(\B_DOUT_TEMPR100[1] ), 
        .C(\B_DOUT_TEMPR101[1] ), .D(\B_DOUT_TEMPR102[1] ), .Y(
        OR4_1151_Y));
    OR4 OR4_682 (.A(\A_DOUT_TEMPR87[18] ), .B(\A_DOUT_TEMPR88[18] ), 
        .C(\A_DOUT_TEMPR89[18] ), .D(\A_DOUT_TEMPR90[18] ), .Y(
        OR4_682_Y));
    OR4 OR4_447 (.A(\B_DOUT_TEMPR20[14] ), .B(\B_DOUT_TEMPR21[14] ), 
        .C(\B_DOUT_TEMPR22[14] ), .D(\B_DOUT_TEMPR23[14] ), .Y(
        OR4_447_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%38%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R38C3 (
        .A_DOUT({nc22890, nc22891, nc22892, nc22893, nc22894, nc22895, 
        nc22896, nc22897, nc22898, nc22899, nc22900, nc22901, nc22902, 
        nc22903, nc22904, \A_DOUT_TEMPR38[19] , \A_DOUT_TEMPR38[18] , 
        \A_DOUT_TEMPR38[17] , \A_DOUT_TEMPR38[16] , 
        \A_DOUT_TEMPR38[15] }), .B_DOUT({nc22905, nc22906, nc22907, 
        nc22908, nc22909, nc22910, nc22911, nc22912, nc22913, nc22914, 
        nc22915, nc22916, nc22917, nc22918, nc22919, 
        \B_DOUT_TEMPR38[19] , \B_DOUT_TEMPR38[18] , 
        \B_DOUT_TEMPR38[17] , \B_DOUT_TEMPR38[16] , 
        \B_DOUT_TEMPR38[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[38][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%84%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R84C4 (
        .A_DOUT({nc22920, nc22921, nc22922, nc22923, nc22924, nc22925, 
        nc22926, nc22927, nc22928, nc22929, nc22930, nc22931, nc22932, 
        nc22933, nc22934, \A_DOUT_TEMPR84[24] , \A_DOUT_TEMPR84[23] , 
        \A_DOUT_TEMPR84[22] , \A_DOUT_TEMPR84[21] , 
        \A_DOUT_TEMPR84[20] }), .B_DOUT({nc22935, nc22936, nc22937, 
        nc22938, nc22939, nc22940, nc22941, nc22942, nc22943, nc22944, 
        nc22945, nc22946, nc22947, nc22948, nc22949, 
        \B_DOUT_TEMPR84[24] , \B_DOUT_TEMPR84[23] , 
        \B_DOUT_TEMPR84[22] , \B_DOUT_TEMPR84[21] , 
        \B_DOUT_TEMPR84[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[84][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1375 (.A(\B_DOUT_TEMPR24[13] ), .B(\B_DOUT_TEMPR25[13] ), 
        .C(\B_DOUT_TEMPR26[13] ), .D(\B_DOUT_TEMPR27[13] ), .Y(
        OR4_1375_Y));
    OR4 OR4_2126 (.A(\A_DOUT_TEMPR75[28] ), .B(\A_DOUT_TEMPR76[28] ), 
        .C(\A_DOUT_TEMPR77[28] ), .D(\A_DOUT_TEMPR78[28] ), .Y(
        OR4_2126_Y));
    OR4 OR4_21 (.A(\A_DOUT_TEMPR79[36] ), .B(\A_DOUT_TEMPR80[36] ), .C(
        \A_DOUT_TEMPR81[36] ), .D(\A_DOUT_TEMPR82[36] ), .Y(OR4_21_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[15]  (.A(CFG3_13_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[15] ));
    OR4 OR4_1443 (.A(\B_DOUT_TEMPR111[34] ), .B(\B_DOUT_TEMPR112[34] ), 
        .C(\B_DOUT_TEMPR113[34] ), .D(\B_DOUT_TEMPR114[34] ), .Y(
        OR4_1443_Y));
    OR4 OR4_1055 (.A(\B_DOUT_TEMPR40[36] ), .B(\B_DOUT_TEMPR41[36] ), 
        .C(\B_DOUT_TEMPR42[36] ), .D(\B_DOUT_TEMPR43[36] ), .Y(
        OR4_1055_Y));
    OR4 OR4_2528 (.A(\A_DOUT_TEMPR103[32] ), .B(\A_DOUT_TEMPR104[32] ), 
        .C(\A_DOUT_TEMPR105[32] ), .D(\A_DOUT_TEMPR106[32] ), .Y(
        OR4_2528_Y));
    OR4 OR4_232 (.A(OR4_26_Y), .B(OR4_832_Y), .C(OR4_2949_Y), .D(
        OR4_2938_Y), .Y(OR4_232_Y));
    OR4 OR4_2877 (.A(\A_DOUT_TEMPR79[16] ), .B(\A_DOUT_TEMPR80[16] ), 
        .C(\A_DOUT_TEMPR81[16] ), .D(\A_DOUT_TEMPR82[16] ), .Y(
        OR4_2877_Y));
    OR4 OR4_1003 (.A(\A_DOUT_TEMPR24[8] ), .B(\A_DOUT_TEMPR25[8] ), .C(
        \A_DOUT_TEMPR26[8] ), .D(\A_DOUT_TEMPR27[8] ), .Y(OR4_1003_Y));
    OR4 OR4_117 (.A(\A_DOUT_TEMPR107[19] ), .B(\A_DOUT_TEMPR108[19] ), 
        .C(\A_DOUT_TEMPR109[19] ), .D(\A_DOUT_TEMPR110[19] ), .Y(
        OR4_117_Y));
    OR4 OR4_1216 (.A(OR4_224_Y), .B(OR4_2450_Y), .C(OR4_1627_Y), .D(
        OR4_571_Y), .Y(OR4_1216_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%34%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R34C1 (
        .A_DOUT({nc22950, nc22951, nc22952, nc22953, nc22954, nc22955, 
        nc22956, nc22957, nc22958, nc22959, nc22960, nc22961, nc22962, 
        nc22963, nc22964, \A_DOUT_TEMPR34[9] , \A_DOUT_TEMPR34[8] , 
        \A_DOUT_TEMPR34[7] , \A_DOUT_TEMPR34[6] , \A_DOUT_TEMPR34[5] })
        , .B_DOUT({nc22965, nc22966, nc22967, nc22968, nc22969, 
        nc22970, nc22971, nc22972, nc22973, nc22974, nc22975, nc22976, 
        nc22977, nc22978, nc22979, \B_DOUT_TEMPR34[9] , 
        \B_DOUT_TEMPR34[8] , \B_DOUT_TEMPR34[7] , \B_DOUT_TEMPR34[6] , 
        \B_DOUT_TEMPR34[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[34][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[5]  (.A(CFG3_1_Y), .B(CFG3_14_Y)
        , .Y(\BLKX2[5] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%30%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R30C4 (
        .A_DOUT({nc22980, nc22981, nc22982, nc22983, nc22984, nc22985, 
        nc22986, nc22987, nc22988, nc22989, nc22990, nc22991, nc22992, 
        nc22993, nc22994, \A_DOUT_TEMPR30[24] , \A_DOUT_TEMPR30[23] , 
        \A_DOUT_TEMPR30[22] , \A_DOUT_TEMPR30[21] , 
        \A_DOUT_TEMPR30[20] }), .B_DOUT({nc22995, nc22996, nc22997, 
        nc22998, nc22999, nc23000, nc23001, nc23002, nc23003, nc23004, 
        nc23005, nc23006, nc23007, nc23008, nc23009, 
        \B_DOUT_TEMPR30[24] , \B_DOUT_TEMPR30[23] , 
        \B_DOUT_TEMPR30[22] , \B_DOUT_TEMPR30[21] , 
        \B_DOUT_TEMPR30[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1601 (.A(OR4_1905_Y), .B(OR4_1252_Y), .C(OR2_2_Y), .D(
        \B_DOUT_TEMPR74[9] ), .Y(OR4_1601_Y));
    OR2 OR2_6 (.A(\A_DOUT_TEMPR72[34] ), .B(\A_DOUT_TEMPR73[34] ), .Y(
        OR2_6_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%91%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R91C2 (
        .A_DOUT({nc23010, nc23011, nc23012, nc23013, nc23014, nc23015, 
        nc23016, nc23017, nc23018, nc23019, nc23020, nc23021, nc23022, 
        nc23023, nc23024, \A_DOUT_TEMPR91[14] , \A_DOUT_TEMPR91[13] , 
        \A_DOUT_TEMPR91[12] , \A_DOUT_TEMPR91[11] , 
        \A_DOUT_TEMPR91[10] }), .B_DOUT({nc23025, nc23026, nc23027, 
        nc23028, nc23029, nc23030, nc23031, nc23032, nc23033, nc23034, 
        nc23035, nc23036, nc23037, nc23038, nc23039, 
        \B_DOUT_TEMPR91[14] , \B_DOUT_TEMPR91[13] , 
        \B_DOUT_TEMPR91[12] , \B_DOUT_TEMPR91[11] , 
        \B_DOUT_TEMPR91[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[91][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[38]  (.A(OR4_817_Y), .B(OR4_1984_Y), .C(OR4_689_Y), 
        .D(OR4_2560_Y), .Y(B_DOUT[38]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%52%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R52C2 (
        .A_DOUT({nc23040, nc23041, nc23042, nc23043, nc23044, nc23045, 
        nc23046, nc23047, nc23048, nc23049, nc23050, nc23051, nc23052, 
        nc23053, nc23054, \A_DOUT_TEMPR52[14] , \A_DOUT_TEMPR52[13] , 
        \A_DOUT_TEMPR52[12] , \A_DOUT_TEMPR52[11] , 
        \A_DOUT_TEMPR52[10] }), .B_DOUT({nc23055, nc23056, nc23057, 
        nc23058, nc23059, nc23060, nc23061, nc23062, nc23063, nc23064, 
        nc23065, nc23066, nc23067, nc23068, nc23069, 
        \B_DOUT_TEMPR52[14] , \B_DOUT_TEMPR52[13] , 
        \B_DOUT_TEMPR52[12] , \B_DOUT_TEMPR52[11] , 
        \B_DOUT_TEMPR52[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[52][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2405 (.A(\B_DOUT_TEMPR115[11] ), .B(\B_DOUT_TEMPR116[11] ), 
        .C(\B_DOUT_TEMPR117[11] ), .D(\B_DOUT_TEMPR118[11] ), .Y(
        OR4_2405_Y));
    OR4 OR4_1703 (.A(\A_DOUT_TEMPR64[38] ), .B(\A_DOUT_TEMPR65[38] ), 
        .C(\A_DOUT_TEMPR66[38] ), .D(\A_DOUT_TEMPR67[38] ), .Y(
        OR4_1703_Y));
    OR4 \OR4_A_DOUT[12]  (.A(OR4_2577_Y), .B(OR4_1155_Y), .C(
        OR4_2085_Y), .D(OR4_1757_Y), .Y(A_DOUT[12]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%108%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R108C1 (
        .A_DOUT({nc23070, nc23071, nc23072, nc23073, nc23074, nc23075, 
        nc23076, nc23077, nc23078, nc23079, nc23080, nc23081, nc23082, 
        nc23083, nc23084, \A_DOUT_TEMPR108[9] , \A_DOUT_TEMPR108[8] , 
        \A_DOUT_TEMPR108[7] , \A_DOUT_TEMPR108[6] , 
        \A_DOUT_TEMPR108[5] }), .B_DOUT({nc23085, nc23086, nc23087, 
        nc23088, nc23089, nc23090, nc23091, nc23092, nc23093, nc23094, 
        nc23095, nc23096, nc23097, nc23098, nc23099, 
        \B_DOUT_TEMPR108[9] , \B_DOUT_TEMPR108[8] , 
        \B_DOUT_TEMPR108[7] , \B_DOUT_TEMPR108[6] , 
        \B_DOUT_TEMPR108[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[108][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_1 (.A(\B_DOUT_TEMPR72[37] ), .B(\B_DOUT_TEMPR73[37] ), .Y(
        OR2_1_Y));
    OR4 OR4_1105 (.A(\B_DOUT_TEMPR16[27] ), .B(\B_DOUT_TEMPR17[27] ), 
        .C(\B_DOUT_TEMPR18[27] ), .D(\B_DOUT_TEMPR19[27] ), .Y(
        OR4_1105_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%62%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R62C0 (
        .A_DOUT({nc23100, nc23101, nc23102, nc23103, nc23104, nc23105, 
        nc23106, nc23107, nc23108, nc23109, nc23110, nc23111, nc23112, 
        nc23113, nc23114, \A_DOUT_TEMPR62[4] , \A_DOUT_TEMPR62[3] , 
        \A_DOUT_TEMPR62[2] , \A_DOUT_TEMPR62[1] , \A_DOUT_TEMPR62[0] })
        , .B_DOUT({nc23115, nc23116, nc23117, nc23118, nc23119, 
        nc23120, nc23121, nc23122, nc23123, nc23124, nc23125, nc23126, 
        nc23127, nc23128, nc23129, \B_DOUT_TEMPR62[4] , 
        \B_DOUT_TEMPR62[3] , \B_DOUT_TEMPR62[2] , \B_DOUT_TEMPR62[1] , 
        \B_DOUT_TEMPR62[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[62][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[7]  (.A(CFG3_13_Y), .B(
        CFG3_14_Y), .Y(\BLKX2[7] ));
    OR4 OR4_1857 (.A(\B_DOUT_TEMPR107[35] ), .B(\B_DOUT_TEMPR108[35] ), 
        .C(\B_DOUT_TEMPR109[35] ), .D(\B_DOUT_TEMPR110[35] ), .Y(
        OR4_1857_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%76%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R76C5 (
        .A_DOUT({nc23130, nc23131, nc23132, nc23133, nc23134, nc23135, 
        nc23136, nc23137, nc23138, nc23139, nc23140, nc23141, nc23142, 
        nc23143, nc23144, \A_DOUT_TEMPR76[29] , \A_DOUT_TEMPR76[28] , 
        \A_DOUT_TEMPR76[27] , \A_DOUT_TEMPR76[26] , 
        \A_DOUT_TEMPR76[25] }), .B_DOUT({nc23145, nc23146, nc23147, 
        nc23148, nc23149, nc23150, nc23151, nc23152, nc23153, nc23154, 
        nc23155, nc23156, nc23157, nc23158, nc23159, 
        \B_DOUT_TEMPR76[29] , \B_DOUT_TEMPR76[28] , 
        \B_DOUT_TEMPR76[27] , \B_DOUT_TEMPR76[26] , 
        \B_DOUT_TEMPR76[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[76][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%79%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R79C5 (
        .A_DOUT({nc23160, nc23161, nc23162, nc23163, nc23164, nc23165, 
        nc23166, nc23167, nc23168, nc23169, nc23170, nc23171, nc23172, 
        nc23173, nc23174, \A_DOUT_TEMPR79[29] , \A_DOUT_TEMPR79[28] , 
        \A_DOUT_TEMPR79[27] , \A_DOUT_TEMPR79[26] , 
        \A_DOUT_TEMPR79[25] }), .B_DOUT({nc23175, nc23176, nc23177, 
        nc23178, nc23179, nc23180, nc23181, nc23182, nc23183, nc23184, 
        nc23185, nc23186, nc23187, nc23188, nc23189, 
        \B_DOUT_TEMPR79[29] , \B_DOUT_TEMPR79[28] , 
        \B_DOUT_TEMPR79[27] , \B_DOUT_TEMPR79[26] , 
        \B_DOUT_TEMPR79[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[79][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_16 (.A(OR4_1601_Y), .B(OR4_916_Y), .C(OR4_80_Y), .D(
        OR4_2058_Y), .Y(OR4_16_Y));
    OR4 OR4_769 (.A(\B_DOUT_TEMPR83[30] ), .B(\B_DOUT_TEMPR84[30] ), 
        .C(\B_DOUT_TEMPR85[30] ), .D(\B_DOUT_TEMPR86[30] ), .Y(
        OR4_769_Y));
    OR4 OR4_1584 (.A(\A_DOUT_TEMPR36[18] ), .B(\A_DOUT_TEMPR37[18] ), 
        .C(\A_DOUT_TEMPR38[18] ), .D(\A_DOUT_TEMPR39[18] ), .Y(
        OR4_1584_Y));
    OR4 OR4_478 (.A(OR4_441_Y), .B(OR4_742_Y), .C(OR4_381_Y), .D(
        OR4_759_Y), .Y(OR4_478_Y));
    OR4 OR4_2636 (.A(\B_DOUT_TEMPR4[22] ), .B(\B_DOUT_TEMPR5[22] ), .C(
        \B_DOUT_TEMPR6[22] ), .D(\B_DOUT_TEMPR7[22] ), .Y(OR4_2636_Y));
    OR4 OR4_2256 (.A(\A_DOUT_TEMPR83[31] ), .B(\A_DOUT_TEMPR84[31] ), 
        .C(\A_DOUT_TEMPR85[31] ), .D(\A_DOUT_TEMPR86[31] ), .Y(
        OR4_2256_Y));
    OR4 OR4_574 (.A(\B_DOUT_TEMPR32[38] ), .B(\B_DOUT_TEMPR33[38] ), 
        .C(\B_DOUT_TEMPR34[38] ), .D(\B_DOUT_TEMPR35[38] ), .Y(
        OR4_574_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%108%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R108C3 (
        .A_DOUT({nc23190, nc23191, nc23192, nc23193, nc23194, nc23195, 
        nc23196, nc23197, nc23198, nc23199, nc23200, nc23201, nc23202, 
        nc23203, nc23204, \A_DOUT_TEMPR108[19] , \A_DOUT_TEMPR108[18] , 
        \A_DOUT_TEMPR108[17] , \A_DOUT_TEMPR108[16] , 
        \A_DOUT_TEMPR108[15] }), .B_DOUT({nc23205, nc23206, nc23207, 
        nc23208, nc23209, nc23210, nc23211, nc23212, nc23213, nc23214, 
        nc23215, nc23216, nc23217, nc23218, nc23219, 
        \B_DOUT_TEMPR108[19] , \B_DOUT_TEMPR108[18] , 
        \B_DOUT_TEMPR108[17] , \B_DOUT_TEMPR108[16] , 
        \B_DOUT_TEMPR108[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[108][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%61%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R61C6 (
        .A_DOUT({nc23220, nc23221, nc23222, nc23223, nc23224, nc23225, 
        nc23226, nc23227, nc23228, nc23229, nc23230, nc23231, nc23232, 
        nc23233, nc23234, \A_DOUT_TEMPR61[34] , \A_DOUT_TEMPR61[33] , 
        \A_DOUT_TEMPR61[32] , \A_DOUT_TEMPR61[31] , 
        \A_DOUT_TEMPR61[30] }), .B_DOUT({nc23235, nc23236, nc23237, 
        nc23238, nc23239, nc23240, nc23241, nc23242, nc23243, nc23244, 
        nc23245, nc23246, nc23247, nc23248, nc23249, 
        \B_DOUT_TEMPR61[34] , \B_DOUT_TEMPR61[33] , 
        \B_DOUT_TEMPR61[32] , \B_DOUT_TEMPR61[31] , 
        \B_DOUT_TEMPR61[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[61][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2130 (.A(OR4_2411_Y), .B(OR4_190_Y), .C(OR4_2284_Y), .D(
        OR4_1319_Y), .Y(OR4_2130_Y));
    OR4 OR4_665 (.A(\A_DOUT_TEMPR48[21] ), .B(\A_DOUT_TEMPR49[21] ), 
        .C(\A_DOUT_TEMPR50[21] ), .D(\A_DOUT_TEMPR51[21] ), .Y(
        OR4_665_Y));
    OR4 OR4_1636 (.A(\A_DOUT_TEMPR24[19] ), .B(\A_DOUT_TEMPR25[19] ), 
        .C(\A_DOUT_TEMPR26[19] ), .D(\A_DOUT_TEMPR27[19] ), .Y(
        OR4_1636_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%53%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R53C1 (
        .A_DOUT({nc23250, nc23251, nc23252, nc23253, nc23254, nc23255, 
        nc23256, nc23257, nc23258, nc23259, nc23260, nc23261, nc23262, 
        nc23263, nc23264, \A_DOUT_TEMPR53[9] , \A_DOUT_TEMPR53[8] , 
        \A_DOUT_TEMPR53[7] , \A_DOUT_TEMPR53[6] , \A_DOUT_TEMPR53[5] })
        , .B_DOUT({nc23265, nc23266, nc23267, nc23268, nc23269, 
        nc23270, nc23271, nc23272, nc23273, nc23274, nc23275, nc23276, 
        nc23277, nc23278, nc23279, \B_DOUT_TEMPR53[9] , 
        \B_DOUT_TEMPR53[8] , \B_DOUT_TEMPR53[7] , \B_DOUT_TEMPR53[6] , 
        \B_DOUT_TEMPR53[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[53][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1001 (.A(\A_DOUT_TEMPR16[19] ), .B(\A_DOUT_TEMPR17[19] ), 
        .C(\A_DOUT_TEMPR18[19] ), .D(\A_DOUT_TEMPR19[19] ), .Y(
        OR4_1001_Y));
    OR4 OR4_2706 (.A(\A_DOUT_TEMPR91[8] ), .B(\A_DOUT_TEMPR92[8] ), .C(
        \A_DOUT_TEMPR93[8] ), .D(\A_DOUT_TEMPR94[8] ), .Y(OR4_2706_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[4]  (.A(CFG3_12_Y), .B(
        CFG3_16_Y), .Y(\BLKY2[4] ));
    OR4 OR4_1130 (.A(\B_DOUT_TEMPR91[22] ), .B(\B_DOUT_TEMPR92[22] ), 
        .C(\B_DOUT_TEMPR93[22] ), .D(\B_DOUT_TEMPR94[22] ), .Y(
        OR4_1130_Y));
    OR4 OR4_269 (.A(\B_DOUT_TEMPR99[25] ), .B(\B_DOUT_TEMPR100[25] ), 
        .C(\B_DOUT_TEMPR101[25] ), .D(\B_DOUT_TEMPR102[25] ), .Y(
        OR4_269_Y));
    OR4 OR4_1816 (.A(OR4_2252_Y), .B(OR4_137_Y), .C(OR4_2863_Y), .D(
        OR4_1305_Y), .Y(OR4_1816_Y));
    OR4 OR4_763 (.A(OR4_220_Y), .B(OR4_2269_Y), .C(OR4_2490_Y), .D(
        OR4_2286_Y), .Y(OR4_763_Y));
    OR4 OR4_2017 (.A(\A_DOUT_TEMPR4[21] ), .B(\A_DOUT_TEMPR5[21] ), .C(
        \A_DOUT_TEMPR6[21] ), .D(\A_DOUT_TEMPR7[21] ), .Y(OR4_2017_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%10%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R10C7 (
        .A_DOUT({nc23280, nc23281, nc23282, nc23283, nc23284, nc23285, 
        nc23286, nc23287, nc23288, nc23289, nc23290, nc23291, nc23292, 
        nc23293, nc23294, \A_DOUT_TEMPR10[39] , \A_DOUT_TEMPR10[38] , 
        \A_DOUT_TEMPR10[37] , \A_DOUT_TEMPR10[36] , 
        \A_DOUT_TEMPR10[35] }), .B_DOUT({nc23295, nc23296, nc23297, 
        nc23298, nc23299, nc23300, nc23301, nc23302, nc23303, nc23304, 
        nc23305, nc23306, nc23307, nc23308, nc23309, 
        \B_DOUT_TEMPR10[39] , \B_DOUT_TEMPR10[38] , 
        \B_DOUT_TEMPR10[37] , \B_DOUT_TEMPR10[36] , 
        \B_DOUT_TEMPR10[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%49%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R49C7 (
        .A_DOUT({nc23310, nc23311, nc23312, nc23313, nc23314, nc23315, 
        nc23316, nc23317, nc23318, nc23319, nc23320, nc23321, nc23322, 
        nc23323, nc23324, \A_DOUT_TEMPR49[39] , \A_DOUT_TEMPR49[38] , 
        \A_DOUT_TEMPR49[37] , \A_DOUT_TEMPR49[36] , 
        \A_DOUT_TEMPR49[35] }), .B_DOUT({nc23325, nc23326, nc23327, 
        nc23328, nc23329, nc23330, nc23331, nc23332, nc23333, nc23334, 
        nc23335, nc23336, nc23337, nc23338, nc23339, 
        \B_DOUT_TEMPR49[39] , \B_DOUT_TEMPR49[38] , 
        \B_DOUT_TEMPR49[37] , \B_DOUT_TEMPR49[36] , 
        \B_DOUT_TEMPR49[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2319 (.A(\A_DOUT_TEMPR111[21] ), .B(\A_DOUT_TEMPR112[21] ), 
        .C(\A_DOUT_TEMPR113[21] ), .D(\A_DOUT_TEMPR114[21] ), .Y(
        OR4_2319_Y));
    OR4 OR4_1526 (.A(OR4_494_Y), .B(OR4_2604_Y), .C(OR4_239_Y), .D(
        OR4_547_Y), .Y(OR4_1526_Y));
    OR4 OR4_2217 (.A(OR4_673_Y), .B(OR4_999_Y), .C(OR4_604_Y), .D(
        OR4_1016_Y), .Y(OR4_2217_Y));
    OR4 OR4_1281 (.A(\B_DOUT_TEMPR48[27] ), .B(\B_DOUT_TEMPR49[27] ), 
        .C(\B_DOUT_TEMPR50[27] ), .D(\B_DOUT_TEMPR51[27] ), .Y(
        OR4_1281_Y));
    OR4 OR4_1727 (.A(OR4_1607_Y), .B(OR4_70_Y), .C(OR4_654_Y), .D(
        OR4_465_Y), .Y(OR4_1727_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%92%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R92C3 (
        .A_DOUT({nc23340, nc23341, nc23342, nc23343, nc23344, nc23345, 
        nc23346, nc23347, nc23348, nc23349, nc23350, nc23351, nc23352, 
        nc23353, nc23354, \A_DOUT_TEMPR92[19] , \A_DOUT_TEMPR92[18] , 
        \A_DOUT_TEMPR92[17] , \A_DOUT_TEMPR92[16] , 
        \A_DOUT_TEMPR92[15] }), .B_DOUT({nc23355, nc23356, nc23357, 
        nc23358, nc23359, nc23360, nc23361, nc23362, nc23363, nc23364, 
        nc23365, nc23366, nc23367, nc23368, nc23369, 
        \B_DOUT_TEMPR92[19] , \B_DOUT_TEMPR92[18] , 
        \B_DOUT_TEMPR92[17] , \B_DOUT_TEMPR92[16] , 
        \B_DOUT_TEMPR92[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[92][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2365 (.A(\A_DOUT_TEMPR79[9] ), .B(\A_DOUT_TEMPR80[9] ), .C(
        \A_DOUT_TEMPR81[9] ), .D(\A_DOUT_TEMPR82[9] ), .Y(OR4_2365_Y));
    OR4 OR4_1521 (.A(\A_DOUT_TEMPR64[16] ), .B(\A_DOUT_TEMPR65[16] ), 
        .C(\A_DOUT_TEMPR66[16] ), .D(\A_DOUT_TEMPR67[16] ), .Y(
        OR4_1521_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%32%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R32C2 (
        .A_DOUT({nc23370, nc23371, nc23372, nc23373, nc23374, nc23375, 
        nc23376, nc23377, nc23378, nc23379, nc23380, nc23381, nc23382, 
        nc23383, nc23384, \A_DOUT_TEMPR32[14] , \A_DOUT_TEMPR32[13] , 
        \A_DOUT_TEMPR32[12] , \A_DOUT_TEMPR32[11] , 
        \A_DOUT_TEMPR32[10] }), .B_DOUT({nc23385, nc23386, nc23387, 
        nc23388, nc23389, nc23390, nc23391, nc23392, nc23393, nc23394, 
        nc23395, nc23396, nc23397, nc23398, nc23399, 
        \B_DOUT_TEMPR32[14] , \B_DOUT_TEMPR32[13] , 
        \B_DOUT_TEMPR32[12] , \B_DOUT_TEMPR32[11] , 
        \B_DOUT_TEMPR32[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[32][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%90%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R90C3 (
        .A_DOUT({nc23400, nc23401, nc23402, nc23403, nc23404, nc23405, 
        nc23406, nc23407, nc23408, nc23409, nc23410, nc23411, nc23412, 
        nc23413, nc23414, \A_DOUT_TEMPR90[19] , \A_DOUT_TEMPR90[18] , 
        \A_DOUT_TEMPR90[17] , \A_DOUT_TEMPR90[16] , 
        \A_DOUT_TEMPR90[15] }), .B_DOUT({nc23415, nc23416, nc23417, 
        nc23418, nc23419, nc23420, nc23421, nc23422, nc23423, nc23424, 
        nc23425, nc23426, nc23427, nc23428, nc23429, 
        \B_DOUT_TEMPR90[19] , \B_DOUT_TEMPR90[18] , 
        \B_DOUT_TEMPR90[17] , \B_DOUT_TEMPR90[16] , 
        \B_DOUT_TEMPR90[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[90][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_268 (.A(\A_DOUT_TEMPR75[10] ), .B(\A_DOUT_TEMPR76[10] ), 
        .C(\A_DOUT_TEMPR77[10] ), .D(\A_DOUT_TEMPR78[10] ), .Y(
        OR4_268_Y));
    OR4 OR4_2524 (.A(OR4_2514_Y), .B(OR4_1733_Y), .C(OR4_172_Y), .D(
        OR4_1736_Y), .Y(OR4_2524_Y));
    OR4 OR4_2910 (.A(\B_DOUT_TEMPR16[0] ), .B(\B_DOUT_TEMPR17[0] ), .C(
        \B_DOUT_TEMPR18[0] ), .D(\B_DOUT_TEMPR19[0] ), .Y(OR4_2910_Y));
    OR4 OR4_216 (.A(\A_DOUT_TEMPR40[2] ), .B(\A_DOUT_TEMPR41[2] ), .C(
        \A_DOUT_TEMPR42[2] ), .D(\A_DOUT_TEMPR43[2] ), .Y(OR4_216_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%68%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R68C2 (
        .A_DOUT({nc23430, nc23431, nc23432, nc23433, nc23434, nc23435, 
        nc23436, nc23437, nc23438, nc23439, nc23440, nc23441, nc23442, 
        nc23443, nc23444, \A_DOUT_TEMPR68[14] , \A_DOUT_TEMPR68[13] , 
        \A_DOUT_TEMPR68[12] , \A_DOUT_TEMPR68[11] , 
        \A_DOUT_TEMPR68[10] }), .B_DOUT({nc23445, nc23446, nc23447, 
        nc23448, nc23449, nc23450, nc23451, nc23452, nc23453, nc23454, 
        nc23455, nc23456, nc23457, nc23458, nc23459, 
        \B_DOUT_TEMPR68[14] , \B_DOUT_TEMPR68[13] , 
        \B_DOUT_TEMPR68[12] , \B_DOUT_TEMPR68[11] , 
        \B_DOUT_TEMPR68[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[68][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2856 (.A(\B_DOUT_TEMPR16[1] ), .B(\B_DOUT_TEMPR17[1] ), .C(
        \B_DOUT_TEMPR18[1] ), .D(\B_DOUT_TEMPR19[1] ), .Y(OR4_2856_Y));
    OR4 OR4_408 (.A(OR4_2361_Y), .B(OR4_834_Y), .C(OR4_1415_Y), .D(
        OR4_1243_Y), .Y(OR4_408_Y));
    OR4 OR4_504 (.A(OR4_1939_Y), .B(OR4_1143_Y), .C(OR4_89_Y), .D(
        OR4_397_Y), .Y(OR4_504_Y));
    OR4 OR4_2593 (.A(OR4_2124_Y), .B(OR4_2845_Y), .C(OR4_481_Y), .D(
        OR4_769_Y), .Y(OR4_2593_Y));
    OR4 OR4_1199 (.A(\B_DOUT_TEMPR64[14] ), .B(\B_DOUT_TEMPR65[14] ), 
        .C(\B_DOUT_TEMPR66[14] ), .D(\B_DOUT_TEMPR67[14] ), .Y(
        OR4_1199_Y));
    OR4 OR4_1710 (.A(\B_DOUT_TEMPR115[16] ), .B(\B_DOUT_TEMPR116[16] ), 
        .C(\B_DOUT_TEMPR117[16] ), .D(\B_DOUT_TEMPR118[16] ), .Y(
        OR4_1710_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%114%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R114C0 (
        .A_DOUT({nc23460, nc23461, nc23462, nc23463, nc23464, nc23465, 
        nc23466, nc23467, nc23468, nc23469, nc23470, nc23471, nc23472, 
        nc23473, nc23474, \A_DOUT_TEMPR114[4] , \A_DOUT_TEMPR114[3] , 
        \A_DOUT_TEMPR114[2] , \A_DOUT_TEMPR114[1] , 
        \A_DOUT_TEMPR114[0] }), .B_DOUT({nc23475, nc23476, nc23477, 
        nc23478, nc23479, nc23480, nc23481, nc23482, nc23483, nc23484, 
        nc23485, nc23486, nc23487, nc23488, nc23489, 
        \B_DOUT_TEMPR114[4] , \B_DOUT_TEMPR114[3] , 
        \B_DOUT_TEMPR114[2] , \B_DOUT_TEMPR114[1] , 
        \B_DOUT_TEMPR114[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[114][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1246 (.A(OR4_1576_Y), .B(OR4_88_Y), .C(OR4_956_Y), .D(
        OR4_3000_Y), .Y(OR4_1246_Y));
    OR4 OR4_2193 (.A(\A_DOUT_TEMPR111[1] ), .B(\A_DOUT_TEMPR112[1] ), 
        .C(\A_DOUT_TEMPR113[1] ), .D(\A_DOUT_TEMPR114[1] ), .Y(
        OR4_2193_Y));
    OR4 OR4_579 (.A(OR4_599_Y), .B(OR4_411_Y), .C(OR4_355_Y), .D(
        OR4_2812_Y), .Y(OR4_579_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%96%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R96C6 (
        .A_DOUT({nc23490, nc23491, nc23492, nc23493, nc23494, nc23495, 
        nc23496, nc23497, nc23498, nc23499, nc23500, nc23501, nc23502, 
        nc23503, nc23504, \A_DOUT_TEMPR96[34] , \A_DOUT_TEMPR96[33] , 
        \A_DOUT_TEMPR96[32] , \A_DOUT_TEMPR96[31] , 
        \A_DOUT_TEMPR96[30] }), .B_DOUT({nc23505, nc23506, nc23507, 
        nc23508, nc23509, nc23510, nc23511, nc23512, nc23513, nc23514, 
        nc23515, nc23516, nc23517, nc23518, nc23519, 
        \B_DOUT_TEMPR96[34] , \B_DOUT_TEMPR96[33] , 
        \B_DOUT_TEMPR96[32] , \B_DOUT_TEMPR96[31] , 
        \B_DOUT_TEMPR96[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[96][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%33%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R33C1 (
        .A_DOUT({nc23520, nc23521, nc23522, nc23523, nc23524, nc23525, 
        nc23526, nc23527, nc23528, nc23529, nc23530, nc23531, nc23532, 
        nc23533, nc23534, \A_DOUT_TEMPR33[9] , \A_DOUT_TEMPR33[8] , 
        \A_DOUT_TEMPR33[7] , \A_DOUT_TEMPR33[6] , \A_DOUT_TEMPR33[5] })
        , .B_DOUT({nc23535, nc23536, nc23537, nc23538, nc23539, 
        nc23540, nc23541, nc23542, nc23543, nc23544, nc23545, nc23546, 
        nc23547, nc23548, nc23549, \B_DOUT_TEMPR33[9] , 
        \B_DOUT_TEMPR33[8] , \B_DOUT_TEMPR33[7] , \B_DOUT_TEMPR33[6] , 
        \B_DOUT_TEMPR33[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[33][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2092 (.A(\A_DOUT_TEMPR28[28] ), .B(\A_DOUT_TEMPR29[28] ), 
        .C(\A_DOUT_TEMPR30[28] ), .D(\A_DOUT_TEMPR31[28] ), .Y(
        OR4_2092_Y));
    OR4 OR4_2712 (.A(\A_DOUT_TEMPR64[9] ), .B(\A_DOUT_TEMPR65[9] ), .C(
        \A_DOUT_TEMPR66[9] ), .D(\A_DOUT_TEMPR67[9] ), .Y(OR4_2712_Y));
    OR4 OR4_1961 (.A(OR4_2474_Y), .B(OR4_2268_Y), .C(OR4_110_Y), .D(
        OR4_1324_Y), .Y(OR4_1961_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%68%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R68C3 (
        .A_DOUT({nc23550, nc23551, nc23552, nc23553, nc23554, nc23555, 
        nc23556, nc23557, nc23558, nc23559, nc23560, nc23561, nc23562, 
        nc23563, nc23564, \A_DOUT_TEMPR68[19] , \A_DOUT_TEMPR68[18] , 
        \A_DOUT_TEMPR68[17] , \A_DOUT_TEMPR68[16] , 
        \A_DOUT_TEMPR68[15] }), .B_DOUT({nc23565, nc23566, nc23567, 
        nc23568, nc23569, nc23570, nc23571, nc23572, nc23573, nc23574, 
        nc23575, nc23576, nc23577, nc23578, nc23579, 
        \B_DOUT_TEMPR68[19] , \B_DOUT_TEMPR68[18] , 
        \B_DOUT_TEMPR68[17] , \B_DOUT_TEMPR68[16] , 
        \B_DOUT_TEMPR68[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[68][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%82%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R82C7 (
        .A_DOUT({nc23580, nc23581, nc23582, nc23583, nc23584, nc23585, 
        nc23586, nc23587, nc23588, nc23589, nc23590, nc23591, nc23592, 
        nc23593, nc23594, \A_DOUT_TEMPR82[39] , \A_DOUT_TEMPR82[38] , 
        \A_DOUT_TEMPR82[37] , \A_DOUT_TEMPR82[36] , 
        \A_DOUT_TEMPR82[35] }), .B_DOUT({nc23595, nc23596, nc23597, 
        nc23598, nc23599, nc23600, nc23601, nc23602, nc23603, nc23604, 
        nc23605, nc23606, nc23607, nc23608, nc23609, 
        \B_DOUT_TEMPR82[39] , \B_DOUT_TEMPR82[38] , 
        \B_DOUT_TEMPR82[37] , \B_DOUT_TEMPR82[36] , 
        \B_DOUT_TEMPR82[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[82][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2741 (.A(\B_DOUT_TEMPR107[9] ), .B(\B_DOUT_TEMPR108[9] ), 
        .C(\B_DOUT_TEMPR109[9] ), .D(\B_DOUT_TEMPR110[9] ), .Y(
        OR4_2741_Y));
    OR4 OR4_2221 (.A(\B_DOUT_TEMPR0[34] ), .B(\B_DOUT_TEMPR1[34] ), .C(
        \B_DOUT_TEMPR2[34] ), .D(\B_DOUT_TEMPR3[34] ), .Y(OR4_2221_Y));
    OR4 OR4_26 (.A(\B_DOUT_TEMPR103[23] ), .B(\B_DOUT_TEMPR104[23] ), 
        .C(\B_DOUT_TEMPR105[23] ), .D(\B_DOUT_TEMPR106[23] ), .Y(
        OR4_26_Y));
    OR4 OR4_3029 (.A(\A_DOUT_TEMPR0[23] ), .B(\A_DOUT_TEMPR1[23] ), .C(
        \A_DOUT_TEMPR2[23] ), .D(\A_DOUT_TEMPR3[23] ), .Y(OR4_3029_Y));
    OR4 OR4_2583 (.A(\B_DOUT_TEMPR79[33] ), .B(\B_DOUT_TEMPR80[33] ), 
        .C(\B_DOUT_TEMPR81[33] ), .D(\B_DOUT_TEMPR82[33] ), .Y(
        OR4_2583_Y));
    OR4 OR4_2933 (.A(\B_DOUT_TEMPR16[39] ), .B(\B_DOUT_TEMPR17[39] ), 
        .C(\B_DOUT_TEMPR18[39] ), .D(\B_DOUT_TEMPR19[39] ), .Y(
        OR4_2933_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%64%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R64C1 (
        .A_DOUT({nc23610, nc23611, nc23612, nc23613, nc23614, nc23615, 
        nc23616, nc23617, nc23618, nc23619, nc23620, nc23621, nc23622, 
        nc23623, nc23624, \A_DOUT_TEMPR64[9] , \A_DOUT_TEMPR64[8] , 
        \A_DOUT_TEMPR64[7] , \A_DOUT_TEMPR64[6] , \A_DOUT_TEMPR64[5] })
        , .B_DOUT({nc23625, nc23626, nc23627, nc23628, nc23629, 
        nc23630, nc23631, nc23632, nc23633, nc23634, nc23635, nc23636, 
        nc23637, nc23638, nc23639, \B_DOUT_TEMPR64[9] , 
        \B_DOUT_TEMPR64[8] , \B_DOUT_TEMPR64[7] , \B_DOUT_TEMPR64[6] , 
        \B_DOUT_TEMPR64[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[64][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_167 (.A(\B_DOUT_TEMPR75[6] ), .B(\B_DOUT_TEMPR76[6] ), .C(
        \B_DOUT_TEMPR77[6] ), .D(\B_DOUT_TEMPR78[6] ), .Y(OR4_167_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%60%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R60C4 (
        .A_DOUT({nc23640, nc23641, nc23642, nc23643, nc23644, nc23645, 
        nc23646, nc23647, nc23648, nc23649, nc23650, nc23651, nc23652, 
        nc23653, nc23654, \A_DOUT_TEMPR60[24] , \A_DOUT_TEMPR60[23] , 
        \A_DOUT_TEMPR60[22] , \A_DOUT_TEMPR60[21] , 
        \A_DOUT_TEMPR60[20] }), .B_DOUT({nc23655, nc23656, nc23657, 
        nc23658, nc23659, nc23660, nc23661, nc23662, nc23663, nc23664, 
        nc23665, nc23666, nc23667, nc23668, nc23669, 
        \B_DOUT_TEMPR60[24] , \B_DOUT_TEMPR60[23] , 
        \B_DOUT_TEMPR60[22] , \B_DOUT_TEMPR60[21] , 
        \B_DOUT_TEMPR60[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[60][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2750 (.A(\B_DOUT_TEMPR12[30] ), .B(\B_DOUT_TEMPR13[30] ), 
        .C(\B_DOUT_TEMPR14[30] ), .D(\B_DOUT_TEMPR15[30] ), .Y(
        OR4_2750_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%104%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R104C3 (
        .A_DOUT({nc23670, nc23671, nc23672, nc23673, nc23674, nc23675, 
        nc23676, nc23677, nc23678, nc23679, nc23680, nc23681, nc23682, 
        nc23683, nc23684, \A_DOUT_TEMPR104[19] , \A_DOUT_TEMPR104[18] , 
        \A_DOUT_TEMPR104[17] , \A_DOUT_TEMPR104[16] , 
        \A_DOUT_TEMPR104[15] }), .B_DOUT({nc23685, nc23686, nc23687, 
        nc23688, nc23689, nc23690, nc23691, nc23692, nc23693, nc23694, 
        nc23695, nc23696, nc23697, nc23698, nc23699, 
        \B_DOUT_TEMPR104[19] , \B_DOUT_TEMPR104[18] , 
        \B_DOUT_TEMPR104[17] , \B_DOUT_TEMPR104[16] , 
        \B_DOUT_TEMPR104[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[104][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2183 (.A(\A_DOUT_TEMPR107[10] ), .B(\A_DOUT_TEMPR108[10] ), 
        .C(\A_DOUT_TEMPR109[10] ), .D(\A_DOUT_TEMPR110[10] ), .Y(
        OR4_2183_Y));
    OR4 OR4_1933 (.A(\B_DOUT_TEMPR83[21] ), .B(\B_DOUT_TEMPR84[21] ), 
        .C(\B_DOUT_TEMPR85[21] ), .D(\B_DOUT_TEMPR86[21] ), .Y(
        OR4_1933_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%7%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R7C5 (
        .A_DOUT({nc23700, nc23701, nc23702, nc23703, nc23704, nc23705, 
        nc23706, nc23707, nc23708, nc23709, nc23710, nc23711, nc23712, 
        nc23713, nc23714, \A_DOUT_TEMPR7[29] , \A_DOUT_TEMPR7[28] , 
        \A_DOUT_TEMPR7[27] , \A_DOUT_TEMPR7[26] , \A_DOUT_TEMPR7[25] })
        , .B_DOUT({nc23715, nc23716, nc23717, nc23718, nc23719, 
        nc23720, nc23721, nc23722, nc23723, nc23724, nc23725, nc23726, 
        nc23727, nc23728, nc23729, \B_DOUT_TEMPR7[29] , 
        \B_DOUT_TEMPR7[28] , \B_DOUT_TEMPR7[27] , \B_DOUT_TEMPR7[26] , 
        \B_DOUT_TEMPR7[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1317 (.A(OR4_1060_Y), .B(OR4_279_Y), .C(OR4_948_Y), .D(
        OR4_99_Y), .Y(OR4_1317_Y));
    OR4 OR4_1212 (.A(\A_DOUT_TEMPR28[9] ), .B(\A_DOUT_TEMPR29[9] ), .C(
        \A_DOUT_TEMPR30[9] ), .D(\A_DOUT_TEMPR31[9] ), .Y(OR4_1212_Y));
    OR4 OR4_2612 (.A(\B_DOUT_TEMPR32[24] ), .B(\B_DOUT_TEMPR33[24] ), 
        .C(\B_DOUT_TEMPR34[24] ), .D(\B_DOUT_TEMPR35[24] ), .Y(
        OR4_2612_Y));
    OR4 OR4_2507 (.A(\B_DOUT_TEMPR95[1] ), .B(\B_DOUT_TEMPR96[1] ), .C(
        \B_DOUT_TEMPR97[1] ), .D(\B_DOUT_TEMPR98[1] ), .Y(OR4_2507_Y));
    OR4 OR4_2082 (.A(\B_DOUT_TEMPR32[1] ), .B(\B_DOUT_TEMPR33[1] ), .C(
        \B_DOUT_TEMPR34[1] ), .D(\B_DOUT_TEMPR35[1] ), .Y(OR4_2082_Y));
    OR4 OR4_52 (.A(OR4_468_Y), .B(OR4_1963_Y), .C(OR4_2544_Y), .D(
        OR4_2350_Y), .Y(OR4_52_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%12%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R12C0 (
        .A_DOUT({nc23730, nc23731, nc23732, nc23733, nc23734, nc23735, 
        nc23736, nc23737, nc23738, nc23739, nc23740, nc23741, nc23742, 
        nc23743, nc23744, \A_DOUT_TEMPR12[4] , \A_DOUT_TEMPR12[3] , 
        \A_DOUT_TEMPR12[2] , \A_DOUT_TEMPR12[1] , \A_DOUT_TEMPR12[0] })
        , .B_DOUT({nc23745, nc23746, nc23747, nc23748, nc23749, 
        nc23750, nc23751, nc23752, nc23753, nc23754, nc23755, nc23756, 
        nc23757, nc23758, nc23759, \B_DOUT_TEMPR12[4] , 
        \B_DOUT_TEMPR12[3] , \B_DOUT_TEMPR12[2] , \B_DOUT_TEMPR12[1] , 
        \B_DOUT_TEMPR12[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2331 (.A(\B_DOUT_TEMPR75[7] ), .B(\B_DOUT_TEMPR76[7] ), .C(
        \B_DOUT_TEMPR77[7] ), .D(\B_DOUT_TEMPR78[7] ), .Y(OR4_2331_Y));
    OR4 OR4_1846 (.A(\B_DOUT_TEMPR91[29] ), .B(\B_DOUT_TEMPR92[29] ), 
        .C(\B_DOUT_TEMPR93[29] ), .D(\B_DOUT_TEMPR94[29] ), .Y(
        OR4_1846_Y));
    OR4 OR4_2912 (.A(\B_DOUT_TEMPR75[35] ), .B(\B_DOUT_TEMPR76[35] ), 
        .C(\B_DOUT_TEMPR77[35] ), .D(\B_DOUT_TEMPR78[35] ), .Y(
        OR4_2912_Y));
    OR4 OR4_1263 (.A(\A_DOUT_TEMPR40[31] ), .B(\A_DOUT_TEMPR41[31] ), 
        .C(\A_DOUT_TEMPR42[31] ), .D(\A_DOUT_TEMPR43[31] ), .Y(
        OR4_1263_Y));
    OR4 OR4_509 (.A(\B_DOUT_TEMPR56[14] ), .B(\B_DOUT_TEMPR57[14] ), 
        .C(\B_DOUT_TEMPR58[14] ), .D(\B_DOUT_TEMPR59[14] ), .Y(
        OR4_509_Y));
    OR4 OR4_2831 (.A(\A_DOUT_TEMPR75[9] ), .B(\A_DOUT_TEMPR76[9] ), .C(
        \A_DOUT_TEMPR77[9] ), .D(\A_DOUT_TEMPR78[9] ), .Y(OR4_2831_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%51%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R51C2 (
        .A_DOUT({nc23760, nc23761, nc23762, nc23763, nc23764, nc23765, 
        nc23766, nc23767, nc23768, nc23769, nc23770, nc23771, nc23772, 
        nc23773, nc23774, \A_DOUT_TEMPR51[14] , \A_DOUT_TEMPR51[13] , 
        \A_DOUT_TEMPR51[12] , \A_DOUT_TEMPR51[11] , 
        \A_DOUT_TEMPR51[10] }), .B_DOUT({nc23775, nc23776, nc23777, 
        nc23778, nc23779, nc23780, nc23781, nc23782, nc23783, nc23784, 
        nc23785, nc23786, nc23787, nc23788, nc23789, 
        \B_DOUT_TEMPR51[14] , \B_DOUT_TEMPR51[13] , 
        \B_DOUT_TEMPR51[12] , \B_DOUT_TEMPR51[11] , 
        \B_DOUT_TEMPR51[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[51][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1331 (.A(\A_DOUT_TEMPR111[16] ), .B(\A_DOUT_TEMPR112[16] ), 
        .C(\A_DOUT_TEMPR113[16] ), .D(\A_DOUT_TEMPR114[16] ), .Y(
        OR4_1331_Y));
    OR4 OR4_919 (.A(\B_DOUT_TEMPR52[32] ), .B(\B_DOUT_TEMPR53[32] ), 
        .C(\B_DOUT_TEMPR54[32] ), .D(\B_DOUT_TEMPR55[32] ), .Y(
        OR4_919_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%11%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R11C6 (
        .A_DOUT({nc23790, nc23791, nc23792, nc23793, nc23794, nc23795, 
        nc23796, nc23797, nc23798, nc23799, nc23800, nc23801, nc23802, 
        nc23803, nc23804, \A_DOUT_TEMPR11[34] , \A_DOUT_TEMPR11[33] , 
        \A_DOUT_TEMPR11[32] , \A_DOUT_TEMPR11[31] , 
        \A_DOUT_TEMPR11[30] }), .B_DOUT({nc23805, nc23806, nc23807, 
        nc23808, nc23809, nc23810, nc23811, nc23812, nc23813, nc23814, 
        nc23815, nc23816, nc23817, nc23818, nc23819, 
        \B_DOUT_TEMPR11[34] , \B_DOUT_TEMPR11[33] , 
        \B_DOUT_TEMPR11[32] , \B_DOUT_TEMPR11[31] , 
        \B_DOUT_TEMPR11[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[6]  (.A(CFG3_0_Y), .B(CFG3_14_Y)
        , .Y(\BLKX2[6] ));
    OR4 OR4_382 (.A(OR4_2925_Y), .B(OR4_933_Y), .C(OR4_2621_Y), .D(
        OR4_1030_Y), .Y(OR4_382_Y));
    OR4 OR4_1831 (.A(\B_DOUT_TEMPR83[22] ), .B(\B_DOUT_TEMPR84[22] ), 
        .C(\B_DOUT_TEMPR85[22] ), .D(\B_DOUT_TEMPR86[22] ), .Y(
        OR4_1831_Y));
    OR4 \OR4_B_DOUT[6]  (.A(OR4_652_Y), .B(OR4_168_Y), .C(OR4_1295_Y), 
        .D(OR4_1259_Y), .Y(B_DOUT[6]));
    OR4 OR4_2443 (.A(OR4_3033_Y), .B(OR4_253_Y), .C(OR4_976_Y), .D(
        OR4_1268_Y), .Y(OR4_2443_Y));
    OR4 OR4_1414 (.A(\B_DOUT_TEMPR40[1] ), .B(\B_DOUT_TEMPR41[1] ), .C(
        \B_DOUT_TEMPR42[1] ), .D(\B_DOUT_TEMPR43[1] ), .Y(OR4_1414_Y));
    OR4 OR4_1573 (.A(\A_DOUT_TEMPR0[31] ), .B(\A_DOUT_TEMPR1[31] ), .C(
        \A_DOUT_TEMPR2[31] ), .D(\A_DOUT_TEMPR3[31] ), .Y(OR4_1573_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%108%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R108C6 (
        .A_DOUT({nc23820, nc23821, nc23822, nc23823, nc23824, nc23825, 
        nc23826, nc23827, nc23828, nc23829, nc23830, nc23831, nc23832, 
        nc23833, nc23834, \A_DOUT_TEMPR108[34] , \A_DOUT_TEMPR108[33] , 
        \A_DOUT_TEMPR108[32] , \A_DOUT_TEMPR108[31] , 
        \A_DOUT_TEMPR108[30] }), .B_DOUT({nc23835, nc23836, nc23837, 
        nc23838, nc23839, nc23840, nc23841, nc23842, nc23843, nc23844, 
        nc23845, nc23846, nc23847, nc23848, nc23849, 
        \B_DOUT_TEMPR108[34] , \B_DOUT_TEMPR108[33] , 
        \B_DOUT_TEMPR108[32] , \B_DOUT_TEMPR108[31] , 
        \B_DOUT_TEMPR108[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[108][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%23%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R23C2 (
        .A_DOUT({nc23850, nc23851, nc23852, nc23853, nc23854, nc23855, 
        nc23856, nc23857, nc23858, nc23859, nc23860, nc23861, nc23862, 
        nc23863, nc23864, \A_DOUT_TEMPR23[14] , \A_DOUT_TEMPR23[13] , 
        \A_DOUT_TEMPR23[12] , \A_DOUT_TEMPR23[11] , 
        \A_DOUT_TEMPR23[10] }), .B_DOUT({nc23865, nc23866, nc23867, 
        nc23868, nc23869, nc23870, nc23871, nc23872, nc23873, nc23874, 
        nc23875, nc23876, nc23877, nc23878, nc23879, 
        \B_DOUT_TEMPR23[14] , \B_DOUT_TEMPR23[13] , 
        \B_DOUT_TEMPR23[12] , \B_DOUT_TEMPR23[11] , 
        \B_DOUT_TEMPR23[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2357 (.A(\A_DOUT_TEMPR20[22] ), .B(\A_DOUT_TEMPR21[22] ), 
        .C(\A_DOUT_TEMPR22[22] ), .D(\A_DOUT_TEMPR23[22] ), .Y(
        OR4_2357_Y));
    OR4 OR4_2252 (.A(\A_DOUT_TEMPR48[35] ), .B(\A_DOUT_TEMPR49[35] ), 
        .C(\A_DOUT_TEMPR50[35] ), .D(\A_DOUT_TEMPR51[35] ), .Y(
        OR4_2252_Y));
    OR4 OR4_1173 (.A(\B_DOUT_TEMPR8[33] ), .B(\B_DOUT_TEMPR9[33] ), .C(
        \B_DOUT_TEMPR10[33] ), .D(\B_DOUT_TEMPR11[33] ), .Y(OR4_1173_Y)
        );
    OR4 \OR4_B_DOUT[16]  (.A(OR4_3013_Y), .B(OR4_1892_Y), .C(
        OR4_2588_Y), .D(OR4_924_Y), .Y(B_DOUT[16]));
    OR4 OR4_458 (.A(\B_DOUT_TEMPR56[36] ), .B(\B_DOUT_TEMPR57[36] ), 
        .C(\B_DOUT_TEMPR58[36] ), .D(\B_DOUT_TEMPR59[36] ), .Y(
        OR4_458_Y));
    OR4 OR4_1892 (.A(OR4_1373_Y), .B(OR4_2857_Y), .C(OR4_1285_Y), .D(
        OR4_2861_Y), .Y(OR4_1892_Y));
    OR4 OR4_31 (.A(\B_DOUT_TEMPR28[37] ), .B(\B_DOUT_TEMPR29[37] ), .C(
        \B_DOUT_TEMPR30[37] ), .D(\B_DOUT_TEMPR31[37] ), .Y(OR4_31_Y));
    OR4 OR4_554 (.A(\A_DOUT_TEMPR36[31] ), .B(\A_DOUT_TEMPR37[31] ), 
        .C(\A_DOUT_TEMPR38[31] ), .D(\A_DOUT_TEMPR39[31] ), .Y(
        OR4_554_Y));
    OR4 OR4_1072 (.A(\A_DOUT_TEMPR91[25] ), .B(\A_DOUT_TEMPR92[25] ), 
        .C(\A_DOUT_TEMPR93[25] ), .D(\A_DOUT_TEMPR94[25] ), .Y(
        OR4_1072_Y));
    OR4 OR4_2172 (.A(\A_DOUT_TEMPR115[21] ), .B(\A_DOUT_TEMPR116[21] ), 
        .C(\A_DOUT_TEMPR117[21] ), .D(\A_DOUT_TEMPR118[21] ), .Y(
        OR4_2172_Y));
    OR2 OR2_37 (.A(\B_DOUT_TEMPR72[6] ), .B(\B_DOUT_TEMPR73[6] ), .Y(
        OR2_37_Y));
    OR4 \OR4_A_DOUT[13]  (.A(OR4_2820_Y), .B(OR4_255_Y), .C(OR4_2495_Y)
        , .D(OR4_296_Y), .Y(A_DOUT[13]));
    OR4 OR4_1740 (.A(OR4_244_Y), .B(OR4_2623_Y), .C(OR2_36_Y), .D(
        \B_DOUT_TEMPR74[5] ), .Y(OR4_1740_Y));
    OR2 OR2_52 (.A(\A_DOUT_TEMPR72[13] ), .B(\A_DOUT_TEMPR73[13] ), .Y(
        OR2_52_Y));
    OR4 OR4_1828 (.A(OR4_2109_Y), .B(OR4_8_Y), .C(OR4_2693_Y), .D(
        OR4_1154_Y), .Y(OR4_1828_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%62%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R62C2 (
        .A_DOUT({nc23880, nc23881, nc23882, nc23883, nc23884, nc23885, 
        nc23886, nc23887, nc23888, nc23889, nc23890, nc23891, nc23892, 
        nc23893, nc23894, \A_DOUT_TEMPR62[14] , \A_DOUT_TEMPR62[13] , 
        \A_DOUT_TEMPR62[12] , \A_DOUT_TEMPR62[11] , 
        \A_DOUT_TEMPR62[10] }), .B_DOUT({nc23895, nc23896, nc23897, 
        nc23898, nc23899, nc23900, nc23901, nc23902, nc23903, nc23904, 
        nc23905, nc23906, nc23907, nc23908, nc23909, 
        \B_DOUT_TEMPR62[14] , \B_DOUT_TEMPR62[13] , 
        \B_DOUT_TEMPR62[12] , \B_DOUT_TEMPR62[11] , 
        \B_DOUT_TEMPR62[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[62][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_A_DOUT[28]  (.A(OR4_2821_Y), .B(OR4_2087_Y), .C(
        OR4_1500_Y), .D(OR4_1935_Y), .Y(A_DOUT[28]));
    OR4 OR4_2454 (.A(\A_DOUT_TEMPR87[26] ), .B(\A_DOUT_TEMPR88[26] ), 
        .C(\A_DOUT_TEMPR89[26] ), .D(\A_DOUT_TEMPR90[26] ), .Y(
        OR4_2454_Y));
    OR4 OR4_585 (.A(OR4_115_Y), .B(OR4_1058_Y), .C(OR4_687_Y), .D(
        OR4_2160_Y), .Y(OR4_585_Y));
    OR4 OR4_936 (.A(\A_DOUT_TEMPR115[19] ), .B(\A_DOUT_TEMPR116[19] ), 
        .C(\A_DOUT_TEMPR117[19] ), .D(\A_DOUT_TEMPR118[19] ), .Y(
        OR4_936_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%18%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R18C2 (
        .A_DOUT({nc23910, nc23911, nc23912, nc23913, nc23914, nc23915, 
        nc23916, nc23917, nc23918, nc23919, nc23920, nc23921, nc23922, 
        nc23923, nc23924, \A_DOUT_TEMPR18[14] , \A_DOUT_TEMPR18[13] , 
        \A_DOUT_TEMPR18[12] , \A_DOUT_TEMPR18[11] , 
        \A_DOUT_TEMPR18[10] }), .B_DOUT({nc23925, nc23926, nc23927, 
        nc23928, nc23929, nc23930, nc23931, nc23932, nc23933, nc23934, 
        nc23935, nc23936, nc23937, nc23938, nc23939, 
        \B_DOUT_TEMPR18[14] , \B_DOUT_TEMPR18[13] , 
        \B_DOUT_TEMPR18[12] , \B_DOUT_TEMPR18[11] , 
        \B_DOUT_TEMPR18[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%9%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R9C6 (
        .A_DOUT({nc23940, nc23941, nc23942, nc23943, nc23944, nc23945, 
        nc23946, nc23947, nc23948, nc23949, nc23950, nc23951, nc23952, 
        nc23953, nc23954, \A_DOUT_TEMPR9[34] , \A_DOUT_TEMPR9[33] , 
        \A_DOUT_TEMPR9[32] , \A_DOUT_TEMPR9[31] , \A_DOUT_TEMPR9[30] })
        , .B_DOUT({nc23955, nc23956, nc23957, nc23958, nc23959, 
        nc23960, nc23961, nc23962, nc23963, nc23964, nc23965, nc23966, 
        nc23967, nc23968, nc23969, \B_DOUT_TEMPR9[34] , 
        \B_DOUT_TEMPR9[33] , \B_DOUT_TEMPR9[32] , \B_DOUT_TEMPR9[31] , 
        \B_DOUT_TEMPR9[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2208 (.A(\A_DOUT_TEMPR16[18] ), .B(\A_DOUT_TEMPR17[18] ), 
        .C(\A_DOUT_TEMPR18[18] ), .D(\A_DOUT_TEMPR19[18] ), .Y(
        OR4_2208_Y));
    OR4 OR4_266 (.A(\B_DOUT_TEMPR60[31] ), .B(\B_DOUT_TEMPR61[31] ), 
        .C(\B_DOUT_TEMPR62[31] ), .D(\B_DOUT_TEMPR63[31] ), .Y(
        OR4_266_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%29%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R29C4 (
        .A_DOUT({nc23970, nc23971, nc23972, nc23973, nc23974, nc23975, 
        nc23976, nc23977, nc23978, nc23979, nc23980, nc23981, nc23982, 
        nc23983, nc23984, \A_DOUT_TEMPR29[24] , \A_DOUT_TEMPR29[23] , 
        \A_DOUT_TEMPR29[22] , \A_DOUT_TEMPR29[21] , 
        \A_DOUT_TEMPR29[20] }), .B_DOUT({nc23985, nc23986, nc23987, 
        nc23988, nc23989, nc23990, nc23991, nc23992, nc23993, nc23994, 
        nc23995, nc23996, nc23997, nc23998, nc23999, 
        \B_DOUT_TEMPR29[24] , \B_DOUT_TEMPR29[23] , 
        \B_DOUT_TEMPR29[22] , \B_DOUT_TEMPR29[21] , 
        \B_DOUT_TEMPR29[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[29][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_54 (.A(\A_DOUT_TEMPR16[9] ), .B(\A_DOUT_TEMPR17[9] ), .C(
        \A_DOUT_TEMPR18[9] ), .D(\A_DOUT_TEMPR19[9] ), .Y(OR4_54_Y));
    OR4 OR4_1152 (.A(OR4_498_Y), .B(OR4_1481_Y), .C(OR4_1082_Y), .D(
        OR4_2759_Y), .Y(OR4_1152_Y));
    OR4 OR4_1693 (.A(OR4_2591_Y), .B(OR4_2900_Y), .C(OR4_1435_Y), .D(
        OR4_2348_Y), .Y(OR4_1693_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%52%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R52C3 (
        .A_DOUT({nc24000, nc24001, nc24002, nc24003, nc24004, nc24005, 
        nc24006, nc24007, nc24008, nc24009, nc24010, nc24011, nc24012, 
        nc24013, nc24014, \A_DOUT_TEMPR52[19] , \A_DOUT_TEMPR52[18] , 
        \A_DOUT_TEMPR52[17] , \A_DOUT_TEMPR52[16] , 
        \A_DOUT_TEMPR52[15] }), .B_DOUT({nc24015, nc24016, nc24017, 
        nc24018, nc24019, nc24020, nc24021, nc24022, nc24023, nc24024, 
        nc24025, nc24026, nc24027, nc24028, nc24029, 
        \B_DOUT_TEMPR52[19] , \B_DOUT_TEMPR52[18] , 
        \B_DOUT_TEMPR52[17] , \B_DOUT_TEMPR52[16] , 
        \B_DOUT_TEMPR52[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[52][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_473 (.A(\B_DOUT_TEMPR75[19] ), .B(\B_DOUT_TEMPR76[19] ), 
        .C(\B_DOUT_TEMPR77[19] ), .D(\B_DOUT_TEMPR78[19] ), .Y(
        OR4_473_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%31%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R31C2 (
        .A_DOUT({nc24030, nc24031, nc24032, nc24033, nc24034, nc24035, 
        nc24036, nc24037, nc24038, nc24039, nc24040, nc24041, nc24042, 
        nc24043, nc24044, \A_DOUT_TEMPR31[14] , \A_DOUT_TEMPR31[13] , 
        \A_DOUT_TEMPR31[12] , \A_DOUT_TEMPR31[11] , 
        \A_DOUT_TEMPR31[10] }), .B_DOUT({nc24045, nc24046, nc24047, 
        nc24048, nc24049, nc24050, nc24051, nc24052, nc24053, nc24054, 
        nc24055, nc24056, nc24057, nc24058, nc24059, 
        \B_DOUT_TEMPR31[14] , \B_DOUT_TEMPR31[13] , 
        \B_DOUT_TEMPR31[12] , \B_DOUT_TEMPR31[11] , 
        \B_DOUT_TEMPR31[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_622 (.A(\B_DOUT_TEMPR0[0] ), .B(\B_DOUT_TEMPR1[0] ), .C(
        \B_DOUT_TEMPR2[0] ), .D(\B_DOUT_TEMPR3[0] ), .Y(OR4_622_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%50%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R50C3 (
        .A_DOUT({nc24060, nc24061, nc24062, nc24063, nc24064, nc24065, 
        nc24066, nc24067, nc24068, nc24069, nc24070, nc24071, nc24072, 
        nc24073, nc24074, \A_DOUT_TEMPR50[19] , \A_DOUT_TEMPR50[18] , 
        \A_DOUT_TEMPR50[17] , \A_DOUT_TEMPR50[16] , 
        \A_DOUT_TEMPR50[15] }), .B_DOUT({nc24075, nc24076, nc24077, 
        nc24078, nc24079, nc24080, nc24081, nc24082, nc24083, nc24084, 
        nc24085, nc24086, nc24087, nc24088, nc24089, 
        \B_DOUT_TEMPR50[19] , \B_DOUT_TEMPR50[18] , 
        \B_DOUT_TEMPR50[17] , \B_DOUT_TEMPR50[16] , 
        \B_DOUT_TEMPR50[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[50][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1999 (.A(\A_DOUT_TEMPR28[37] ), .B(\A_DOUT_TEMPR29[37] ), 
        .C(\A_DOUT_TEMPR30[37] ), .D(\A_DOUT_TEMPR31[37] ), .Y(
        OR4_1999_Y));
    OR4 OR4_2419 (.A(OR4_1600_Y), .B(OR4_632_Y), .C(OR4_841_Y), .D(
        OR4_643_Y), .Y(OR4_2419_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENB[12]  (.A(B_WBYTE_EN[6]), .B(
        B_WEN), .Y(\WBYTEENB[12] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%63%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R63C1 (
        .A_DOUT({nc24090, nc24091, nc24092, nc24093, nc24094, nc24095, 
        nc24096, nc24097, nc24098, nc24099, nc24100, nc24101, nc24102, 
        nc24103, nc24104, \A_DOUT_TEMPR63[9] , \A_DOUT_TEMPR63[8] , 
        \A_DOUT_TEMPR63[7] , \A_DOUT_TEMPR63[6] , \A_DOUT_TEMPR63[5] })
        , .B_DOUT({nc24105, nc24106, nc24107, nc24108, nc24109, 
        nc24110, nc24111, nc24112, nc24113, nc24114, nc24115, nc24116, 
        nc24117, nc24118, nc24119, \B_DOUT_TEMPR63[9] , 
        \B_DOUT_TEMPR63[8] , \B_DOUT_TEMPR63[7] , \B_DOUT_TEMPR63[6] , 
        \B_DOUT_TEMPR63[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[63][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1605 (.A(\A_DOUT_TEMPR111[23] ), .B(\A_DOUT_TEMPR112[23] ), 
        .C(\A_DOUT_TEMPR113[23] ), .D(\A_DOUT_TEMPR114[23] ), .Y(
        OR4_1605_Y));
    OR4 OR4_1214 (.A(OR4_1900_Y), .B(OR4_165_Y), .C(OR4_2883_Y), .D(
        OR4_893_Y), .Y(OR4_1214_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%18%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R18C3 (
        .A_DOUT({nc24120, nc24121, nc24122, nc24123, nc24124, nc24125, 
        nc24126, nc24127, nc24128, nc24129, nc24130, nc24131, nc24132, 
        nc24133, nc24134, \A_DOUT_TEMPR18[19] , \A_DOUT_TEMPR18[18] , 
        \A_DOUT_TEMPR18[17] , \A_DOUT_TEMPR18[16] , 
        \A_DOUT_TEMPR18[15] }), .B_DOUT({nc24135, nc24136, nc24137, 
        nc24138, nc24139, nc24140, nc24141, nc24142, nc24143, nc24144, 
        nc24145, nc24146, nc24147, nc24148, nc24149, 
        \B_DOUT_TEMPR18[19] , \B_DOUT_TEMPR18[18] , 
        \B_DOUT_TEMPR18[17] , \B_DOUT_TEMPR18[16] , 
        \B_DOUT_TEMPR18[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[18][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1347 (.A(OR4_1308_Y), .B(OR4_303_Y), .C(OR4_528_Y), .D(
        OR4_322_Y), .Y(OR4_1347_Y));
    OR4 OR4_1242 (.A(\B_DOUT_TEMPR32[10] ), .B(\B_DOUT_TEMPR33[10] ), 
        .C(\B_DOUT_TEMPR34[10] ), .D(\B_DOUT_TEMPR35[10] ), .Y(
        OR4_1242_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_13 (.A(A_ADDR[16]), .B(A_ADDR[15]), 
        .C(A_ADDR[14]), .Y(CFG3_13_Y));
    OR2 OR2_30 (.A(\A_DOUT_TEMPR72[17] ), .B(\A_DOUT_TEMPR73[17] ), .Y(
        OR2_30_Y));
    OR4 OR4_2398 (.A(\B_DOUT_TEMPR99[31] ), .B(\B_DOUT_TEMPR100[31] ), 
        .C(\B_DOUT_TEMPR101[31] ), .D(\B_DOUT_TEMPR102[31] ), .Y(
        OR4_2398_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%14%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R14C1 (
        .A_DOUT({nc24150, nc24151, nc24152, nc24153, nc24154, nc24155, 
        nc24156, nc24157, nc24158, nc24159, nc24160, nc24161, nc24162, 
        nc24163, nc24164, \A_DOUT_TEMPR14[9] , \A_DOUT_TEMPR14[8] , 
        \A_DOUT_TEMPR14[7] , \A_DOUT_TEMPR14[6] , \A_DOUT_TEMPR14[5] })
        , .B_DOUT({nc24165, nc24166, nc24167, nc24168, nc24169, 
        nc24170, nc24171, nc24172, nc24173, nc24174, nc24175, nc24176, 
        nc24177, nc24178, nc24179, \B_DOUT_TEMPR14[9] , 
        \B_DOUT_TEMPR14[8] , \B_DOUT_TEMPR14[7] , \B_DOUT_TEMPR14[6] , 
        \B_DOUT_TEMPR14[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%10%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R10C4 (
        .A_DOUT({nc24180, nc24181, nc24182, nc24183, nc24184, nc24185, 
        nc24186, nc24187, nc24188, nc24189, nc24190, nc24191, nc24192, 
        nc24193, nc24194, \A_DOUT_TEMPR10[24] , \A_DOUT_TEMPR10[23] , 
        \A_DOUT_TEMPR10[22] , \A_DOUT_TEMPR10[21] , 
        \A_DOUT_TEMPR10[20] }), .B_DOUT({nc24195, nc24196, nc24197, 
        nc24198, nc24199, nc24200, nc24201, nc24202, nc24203, nc24204, 
        nc24205, nc24206, nc24207, nc24208, nc24209, 
        \B_DOUT_TEMPR10[24] , \B_DOUT_TEMPR10[23] , 
        \B_DOUT_TEMPR10[22] , \B_DOUT_TEMPR10[21] , 
        \B_DOUT_TEMPR10[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%56%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R56C6 (
        .A_DOUT({nc24210, nc24211, nc24212, nc24213, nc24214, nc24215, 
        nc24216, nc24217, nc24218, nc24219, nc24220, nc24221, nc24222, 
        nc24223, nc24224, \A_DOUT_TEMPR56[34] , \A_DOUT_TEMPR56[33] , 
        \A_DOUT_TEMPR56[32] , \A_DOUT_TEMPR56[31] , 
        \A_DOUT_TEMPR56[30] }), .B_DOUT({nc24225, nc24226, nc24227, 
        nc24228, nc24229, nc24230, nc24231, nc24232, nc24233, nc24234, 
        nc24235, nc24236, nc24237, nc24238, nc24239, 
        \B_DOUT_TEMPR56[34] , \B_DOUT_TEMPR56[33] , 
        \B_DOUT_TEMPR56[32] , \B_DOUT_TEMPR56[31] , 
        \B_DOUT_TEMPR56[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[56][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_559 (.A(\B_DOUT_TEMPR68[2] ), .B(\B_DOUT_TEMPR69[2] ), .C(
        \B_DOUT_TEMPR70[2] ), .D(\B_DOUT_TEMPR71[2] ), .Y(OR4_559_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%0%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R0C4 (
        .A_DOUT({nc24240, nc24241, nc24242, nc24243, nc24244, nc24245, 
        nc24246, nc24247, nc24248, nc24249, nc24250, nc24251, nc24252, 
        nc24253, nc24254, \A_DOUT_TEMPR0[24] , \A_DOUT_TEMPR0[23] , 
        \A_DOUT_TEMPR0[22] , \A_DOUT_TEMPR0[21] , \A_DOUT_TEMPR0[20] })
        , .B_DOUT({nc24255, nc24256, nc24257, nc24258, nc24259, 
        nc24260, nc24261, nc24262, nc24263, nc24264, nc24265, nc24266, 
        nc24267, nc24268, nc24269, \B_DOUT_TEMPR0[24] , 
        \B_DOUT_TEMPR0[23] , \B_DOUT_TEMPR0[22] , \B_DOUT_TEMPR0[21] , 
        \B_DOUT_TEMPR0[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2563 (.A(\A_DOUT_TEMPR79[2] ), .B(\A_DOUT_TEMPR80[2] ), .C(
        \A_DOUT_TEMPR81[2] ), .D(\A_DOUT_TEMPR82[2] ), .Y(OR4_2563_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%79%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R79C7 (
        .A_DOUT({nc24270, nc24271, nc24272, nc24273, nc24274, nc24275, 
        nc24276, nc24277, nc24278, nc24279, nc24280, nc24281, nc24282, 
        nc24283, nc24284, \A_DOUT_TEMPR79[39] , \A_DOUT_TEMPR79[38] , 
        \A_DOUT_TEMPR79[37] , \A_DOUT_TEMPR79[36] , 
        \A_DOUT_TEMPR79[35] }), .B_DOUT({nc24285, nc24286, nc24287, 
        nc24288, nc24289, nc24290, nc24291, nc24292, nc24293, nc24294, 
        nc24295, nc24296, nc24297, nc24298, nc24299, 
        \B_DOUT_TEMPR79[39] , \B_DOUT_TEMPR79[38] , 
        \B_DOUT_TEMPR79[37] , \B_DOUT_TEMPR79[36] , 
        \B_DOUT_TEMPR79[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[79][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1794 (.A(OR4_2091_Y), .B(OR4_1895_Y), .C(OR4_2792_Y), .D(
        OR4_944_Y), .Y(OR4_1794_Y));
    OR4 OR4_1728 (.A(\B_DOUT_TEMPR111[30] ), .B(\B_DOUT_TEMPR112[30] ), 
        .C(\B_DOUT_TEMPR113[30] ), .D(\B_DOUT_TEMPR114[30] ), .Y(
        OR4_1728_Y));
    OR4 OR4_1013 (.A(OR4_2409_Y), .B(OR4_185_Y), .C(OR4_2281_Y), .D(
        OR4_1802_Y), .Y(OR4_1013_Y));
    OR4 OR4_2310 (.A(\B_DOUT_TEMPR68[26] ), .B(\B_DOUT_TEMPR69[26] ), 
        .C(\B_DOUT_TEMPR70[26] ), .D(\B_DOUT_TEMPR71[26] ), .Y(
        OR4_2310_Y));
    OR4 OR4_2417 (.A(\B_DOUT_TEMPR99[18] ), .B(\B_DOUT_TEMPR100[18] ), 
        .C(\B_DOUT_TEMPR101[18] ), .D(\B_DOUT_TEMPR102[18] ), .Y(
        OR4_2417_Y));
    OR4 OR4_81 (.A(OR4_1272_Y), .B(OR4_2301_Y), .C(OR4_1003_Y), .D(
        OR4_2394_Y), .Y(OR4_81_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%96%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R96C0 (
        .A_DOUT({nc24300, nc24301, nc24302, nc24303, nc24304, nc24305, 
        nc24306, nc24307, nc24308, nc24309, nc24310, nc24311, nc24312, 
        nc24313, nc24314, \A_DOUT_TEMPR96[4] , \A_DOUT_TEMPR96[3] , 
        \A_DOUT_TEMPR96[2] , \A_DOUT_TEMPR96[1] , \A_DOUT_TEMPR96[0] })
        , .B_DOUT({nc24315, nc24316, nc24317, nc24318, nc24319, 
        nc24320, nc24321, nc24322, nc24323, nc24324, nc24325, nc24326, 
        nc24327, nc24328, nc24329, \B_DOUT_TEMPR96[4] , 
        \B_DOUT_TEMPR96[3] , \B_DOUT_TEMPR96[2] , \B_DOUT_TEMPR96[1] , 
        \B_DOUT_TEMPR96[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[96][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1607 (.A(\B_DOUT_TEMPR16[32] ), .B(\B_DOUT_TEMPR17[32] ), 
        .C(\B_DOUT_TEMPR18[32] ), .D(\B_DOUT_TEMPR19[32] ), .Y(
        OR4_1607_Y));
    OR4 OR4_1491 (.A(OR4_217_Y), .B(OR4_1705_Y), .C(OR4_2289_Y), .D(
        OR4_2106_Y), .Y(OR4_1491_Y));
    OR4 OR4_1611 (.A(OR4_1059_Y), .B(OR4_861_Y), .C(OR4_793_Y), .D(
        OR4_1591_Y), .Y(OR4_1611_Y));
    OR4 OR4_2163 (.A(OR4_2311_Y), .B(OR4_483_Y), .C(OR2_38_Y), .D(
        \A_DOUT_TEMPR74[18] ), .Y(OR4_2163_Y));
    OR2 OR2_54 (.A(\B_DOUT_TEMPR72[38] ), .B(\B_DOUT_TEMPR73[38] ), .Y(
        OR2_54_Y));
    OR4 OR4_1444 (.A(\B_DOUT_TEMPR107[18] ), .B(\B_DOUT_TEMPR108[18] ), 
        .C(\B_DOUT_TEMPR109[18] ), .D(\B_DOUT_TEMPR110[18] ), .Y(
        OR4_1444_Y));
    OR4 OR4_2254 (.A(\B_DOUT_TEMPR12[11] ), .B(\B_DOUT_TEMPR13[11] ), 
        .C(\B_DOUT_TEMPR14[11] ), .D(\B_DOUT_TEMPR15[11] ), .Y(
        OR4_2254_Y));
    OR4 OR4_1713 (.A(OR4_1002_Y), .B(OR4_2652_Y), .C(OR4_2024_Y), .D(
        OR4_1363_Y), .Y(OR4_1713_Y));
    OR4 OR4_2246 (.A(\B_DOUT_TEMPR103[37] ), .B(\B_DOUT_TEMPR104[37] ), 
        .C(\B_DOUT_TEMPR105[37] ), .D(\B_DOUT_TEMPR106[37] ), .Y(
        OR4_2246_Y));
    OR4 OR4_2062 (.A(\A_DOUT_TEMPR32[38] ), .B(\A_DOUT_TEMPR33[38] ), 
        .C(\A_DOUT_TEMPR34[38] ), .D(\A_DOUT_TEMPR35[38] ), .Y(
        OR4_2062_Y));
    OR4 OR4_403 (.A(\A_DOUT_TEMPR103[37] ), .B(\A_DOUT_TEMPR104[37] ), 
        .C(\A_DOUT_TEMPR105[37] ), .D(\A_DOUT_TEMPR106[37] ), .Y(
        OR4_403_Y));
    OR4 OR4_2388 (.A(\B_DOUT_TEMPR48[7] ), .B(\B_DOUT_TEMPR49[7] ), .C(
        \B_DOUT_TEMPR50[7] ), .D(\B_DOUT_TEMPR51[7] ), .Y(OR4_2388_Y));
    OR4 OR4_1115 (.A(OR4_28_Y), .B(OR4_173_Y), .C(OR4_1658_Y), .D(
        OR4_176_Y), .Y(OR4_1115_Y));
    OR4 OR4_2937 (.A(\B_DOUT_TEMPR4[2] ), .B(\B_DOUT_TEMPR5[2] ), .C(
        \B_DOUT_TEMPR6[2] ), .D(\B_DOUT_TEMPR7[2] ), .Y(OR4_2937_Y));
    OR4 \OR4_A_DOUT[27]  (.A(OR4_180_Y), .B(OR4_1971_Y), .C(OR4_977_Y), 
        .D(OR4_2130_Y), .Y(A_DOUT[27]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%107%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R107C3 (
        .A_DOUT({nc24330, nc24331, nc24332, nc24333, nc24334, nc24335, 
        nc24336, nc24337, nc24338, nc24339, nc24340, nc24341, nc24342, 
        nc24343, nc24344, \A_DOUT_TEMPR107[19] , \A_DOUT_TEMPR107[18] , 
        \A_DOUT_TEMPR107[17] , \A_DOUT_TEMPR107[16] , 
        \A_DOUT_TEMPR107[15] }), .B_DOUT({nc24345, nc24346, nc24347, 
        nc24348, nc24349, nc24350, nc24351, nc24352, nc24353, nc24354, 
        nc24355, nc24356, nc24357, nc24358, nc24359, 
        \B_DOUT_TEMPR107[19] , \B_DOUT_TEMPR107[18] , 
        \B_DOUT_TEMPR107[17] , \B_DOUT_TEMPR107[16] , 
        \B_DOUT_TEMPR107[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[107][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[1]  (.A(CFG3_5_Y), .B(CFG3_14_Y)
        , .Y(\BLKX2[1] ));
    OR4 OR4_969 (.A(OR4_259_Y), .B(OR4_235_Y), .C(OR4_895_Y), .D(
        OR4_63_Y), .Y(OR4_969_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%32%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R32C3 (
        .A_DOUT({nc24360, nc24361, nc24362, nc24363, nc24364, nc24365, 
        nc24366, nc24367, nc24368, nc24369, nc24370, nc24371, nc24372, 
        nc24373, nc24374, \A_DOUT_TEMPR32[19] , \A_DOUT_TEMPR32[18] , 
        \A_DOUT_TEMPR32[17] , \A_DOUT_TEMPR32[16] , 
        \A_DOUT_TEMPR32[15] }), .B_DOUT({nc24375, nc24376, nc24377, 
        nc24378, nc24379, nc24380, nc24381, nc24382, nc24383, nc24384, 
        nc24385, nc24386, nc24387, nc24388, nc24389, 
        \B_DOUT_TEMPR32[19] , \B_DOUT_TEMPR32[18] , 
        \B_DOUT_TEMPR32[17] , \B_DOUT_TEMPR32[16] , 
        \B_DOUT_TEMPR32[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[32][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1937 (.A(\B_DOUT_TEMPR0[6] ), .B(\B_DOUT_TEMPR1[6] ), .C(
        \B_DOUT_TEMPR2[6] ), .D(\B_DOUT_TEMPR3[6] ), .Y(OR4_1937_Y));
    OR4 OR4_498 (.A(\A_DOUT_TEMPR32[7] ), .B(\A_DOUT_TEMPR33[7] ), .C(
        \A_DOUT_TEMPR34[7] ), .D(\A_DOUT_TEMPR35[7] ), .Y(OR4_498_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%30%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R30C3 (
        .A_DOUT({nc24390, nc24391, nc24392, nc24393, nc24394, nc24395, 
        nc24396, nc24397, nc24398, nc24399, nc24400, nc24401, nc24402, 
        nc24403, nc24404, \A_DOUT_TEMPR30[19] , \A_DOUT_TEMPR30[18] , 
        \A_DOUT_TEMPR30[17] , \A_DOUT_TEMPR30[16] , 
        \A_DOUT_TEMPR30[15] }), .B_DOUT({nc24405, nc24406, nc24407, 
        nc24408, nc24409, nc24410, nc24411, nc24412, nc24413, nc24414, 
        nc24415, nc24416, nc24417, nc24418, nc24419, 
        \B_DOUT_TEMPR30[19] , \B_DOUT_TEMPR30[18] , 
        \B_DOUT_TEMPR30[17] , \B_DOUT_TEMPR30[16] , 
        \B_DOUT_TEMPR30[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[30][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2279 (.A(\B_DOUT_TEMPR44[27] ), .B(\B_DOUT_TEMPR45[27] ), 
        .C(\B_DOUT_TEMPR46[27] ), .D(\B_DOUT_TEMPR47[27] ), .Y(
        OR4_2279_Y));
    OR4 OR4_2053 (.A(\A_DOUT_TEMPR0[28] ), .B(\A_DOUT_TEMPR1[28] ), .C(
        \A_DOUT_TEMPR2[28] ), .D(\A_DOUT_TEMPR3[28] ), .Y(OR4_2053_Y));
    OR4 OR4_642 (.A(OR4_921_Y), .B(OR4_1230_Y), .C(OR4_846_Y), .D(
        OR4_1244_Y), .Y(OR4_642_Y));
    OR4 OR4_594 (.A(\B_DOUT_TEMPR64[39] ), .B(\B_DOUT_TEMPR65[39] ), 
        .C(\B_DOUT_TEMPR66[39] ), .D(\B_DOUT_TEMPR67[39] ), .Y(
        OR4_594_Y));
    OR4 OR4_2651 (.A(\A_DOUT_TEMPR16[15] ), .B(\A_DOUT_TEMPR17[15] ), 
        .C(\A_DOUT_TEMPR18[15] ), .D(\A_DOUT_TEMPR19[15] ), .Y(
        OR4_2651_Y));
    OR4 OR4_1011 (.A(\A_DOUT_TEMPR44[22] ), .B(\A_DOUT_TEMPR45[22] ), 
        .C(\A_DOUT_TEMPR46[22] ), .D(\A_DOUT_TEMPR47[22] ), .Y(
        OR4_1011_Y));
    OR4 OR4_1994 (.A(\A_DOUT_TEMPR24[2] ), .B(\A_DOUT_TEMPR25[2] ), .C(
        \A_DOUT_TEMPR26[2] ), .D(\A_DOUT_TEMPR27[2] ), .Y(OR4_1994_Y));
    OR4 OR4_2495 (.A(OR4_420_Y), .B(OR4_2481_Y), .C(OR4_2714_Y), .D(
        OR4_2502_Y), .Y(OR4_2495_Y));
    OR4 OR4_432 (.A(\B_DOUT_TEMPR36[14] ), .B(\B_DOUT_TEMPR37[14] ), 
        .C(\B_DOUT_TEMPR38[14] ), .D(\B_DOUT_TEMPR39[14] ), .Y(
        OR4_432_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[3]  (.A(CFG3_23_Y), .B(
        CFG3_14_Y), .Y(\BLKX2[3] ));
    OR4 OR4_2753 (.A(\A_DOUT_TEMPR64[0] ), .B(\A_DOUT_TEMPR65[0] ), .C(
        \A_DOUT_TEMPR66[0] ), .D(\A_DOUT_TEMPR67[0] ), .Y(OR4_2753_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%46%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R46C1 (
        .A_DOUT({nc24420, nc24421, nc24422, nc24423, nc24424, nc24425, 
        nc24426, nc24427, nc24428, nc24429, nc24430, nc24431, nc24432, 
        nc24433, nc24434, \A_DOUT_TEMPR46[9] , \A_DOUT_TEMPR46[8] , 
        \A_DOUT_TEMPR46[7] , \A_DOUT_TEMPR46[6] , \A_DOUT_TEMPR46[5] })
        , .B_DOUT({nc24435, nc24436, nc24437, nc24438, nc24439, 
        nc24440, nc24441, nc24442, nc24443, nc24444, nc24445, nc24446, 
        nc24447, nc24448, nc24449, \B_DOUT_TEMPR46[9] , 
        \B_DOUT_TEMPR46[8] , \B_DOUT_TEMPR46[7] , \B_DOUT_TEMPR46[6] , 
        \B_DOUT_TEMPR46[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[46][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2830 (.A(OR4_1769_Y), .B(OR4_2982_Y), .C(OR2_30_Y), .D(
        \A_DOUT_TEMPR74[17] ), .Y(OR4_2830_Y));
    OR4 OR4_1996 (.A(\B_DOUT_TEMPR52[4] ), .B(\B_DOUT_TEMPR53[4] ), .C(
        \B_DOUT_TEMPR54[4] ), .D(\B_DOUT_TEMPR55[4] ), .Y(OR4_1996_Y));
    OR4 OR4_36 (.A(\A_DOUT_TEMPR91[34] ), .B(\A_DOUT_TEMPR92[34] ), .C(
        \A_DOUT_TEMPR93[34] ), .D(\A_DOUT_TEMPR94[34] ), .Y(OR4_36_Y));
    OR4 OR4_2155 (.A(\A_DOUT_TEMPR115[18] ), .B(\A_DOUT_TEMPR116[18] ), 
        .C(\A_DOUT_TEMPR117[18] ), .D(\A_DOUT_TEMPR118[18] ), .Y(
        OR4_2155_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%36%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R36C6 (
        .A_DOUT({nc24450, nc24451, nc24452, nc24453, nc24454, nc24455, 
        nc24456, nc24457, nc24458, nc24459, nc24460, nc24461, nc24462, 
        nc24463, nc24464, \A_DOUT_TEMPR36[34] , \A_DOUT_TEMPR36[33] , 
        \A_DOUT_TEMPR36[32] , \A_DOUT_TEMPR36[31] , 
        \A_DOUT_TEMPR36[30] }), .B_DOUT({nc24465, nc24466, nc24467, 
        nc24468, nc24469, nc24470, nc24471, nc24472, nc24473, nc24474, 
        nc24475, nc24476, nc24477, nc24478, nc24479, 
        \B_DOUT_TEMPR36[34] , \B_DOUT_TEMPR36[33] , 
        \B_DOUT_TEMPR36[32] , \B_DOUT_TEMPR36[31] , 
        \B_DOUT_TEMPR36[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1259 (.A(OR4_2685_Y), .B(OR4_1997_Y), .C(OR4_894_Y), .D(
        OR4_2779_Y), .Y(OR4_1259_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%94%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R94C2 (
        .A_DOUT({nc24480, nc24481, nc24482, nc24483, nc24484, nc24485, 
        nc24486, nc24487, nc24488, nc24489, nc24490, nc24491, nc24492, 
        nc24493, nc24494, \A_DOUT_TEMPR94[14] , \A_DOUT_TEMPR94[13] , 
        \A_DOUT_TEMPR94[12] , \A_DOUT_TEMPR94[11] , 
        \A_DOUT_TEMPR94[10] }), .B_DOUT({nc24495, nc24496, nc24497, 
        nc24498, nc24499, nc24500, nc24501, nc24502, nc24503, nc24504, 
        nc24505, nc24506, nc24507, nc24508, nc24509, 
        \B_DOUT_TEMPR94[14] , \B_DOUT_TEMPR94[13] , 
        \B_DOUT_TEMPR94[12] , \B_DOUT_TEMPR94[11] , 
        \B_DOUT_TEMPR94[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[94][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[5]  (.A(CFG3_6_Y), .B(CFG3_16_Y)
        , .Y(\BLKY2[5] ));
    OR4 OR4_2846 (.A(\B_DOUT_TEMPR20[6] ), .B(\B_DOUT_TEMPR21[6] ), .C(
        \B_DOUT_TEMPR22[6] ), .D(\B_DOUT_TEMPR23[6] ), .Y(OR4_2846_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%88%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R88C1 (
        .A_DOUT({nc24510, nc24511, nc24512, nc24513, nc24514, nc24515, 
        nc24516, nc24517, nc24518, nc24519, nc24520, nc24521, nc24522, 
        nc24523, nc24524, \A_DOUT_TEMPR88[9] , \A_DOUT_TEMPR88[8] , 
        \A_DOUT_TEMPR88[7] , \A_DOUT_TEMPR88[6] , \A_DOUT_TEMPR88[5] })
        , .B_DOUT({nc24525, nc24526, nc24527, nc24528, nc24529, 
        nc24530, nc24531, nc24532, nc24533, nc24534, nc24535, nc24536, 
        nc24537, nc24538, nc24539, \B_DOUT_TEMPR88[9] , 
        \B_DOUT_TEMPR88[8] , \B_DOUT_TEMPR88[7] , \B_DOUT_TEMPR88[6] , 
        \B_DOUT_TEMPR88[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[88][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1830 (.A(OR4_428_Y), .B(OR4_729_Y), .C(OR4_369_Y), .D(
        OR4_750_Y), .Y(OR4_1830_Y));
    OR4 OR4_1378 (.A(\A_DOUT_TEMPR87[8] ), .B(\A_DOUT_TEMPR88[8] ), .C(
        \A_DOUT_TEMPR89[8] ), .D(\A_DOUT_TEMPR90[8] ), .Y(OR4_1378_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%12%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R12C2 (
        .A_DOUT({nc24540, nc24541, nc24542, nc24543, nc24544, nc24545, 
        nc24546, nc24547, nc24548, nc24549, nc24550, nc24551, nc24552, 
        nc24553, nc24554, \A_DOUT_TEMPR12[14] , \A_DOUT_TEMPR12[13] , 
        \A_DOUT_TEMPR12[12] , \A_DOUT_TEMPR12[11] , 
        \A_DOUT_TEMPR12[10] }), .B_DOUT({nc24555, nc24556, nc24557, 
        nc24558, nc24559, nc24560, nc24561, nc24562, nc24563, nc24564, 
        nc24565, nc24566, nc24567, nc24568, nc24569, 
        \B_DOUT_TEMPR12[14] , \B_DOUT_TEMPR12[13] , 
        \B_DOUT_TEMPR12[12] , \B_DOUT_TEMPR12[11] , 
        \B_DOUT_TEMPR12[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1761 (.A(OR4_347_Y), .B(OR4_2071_Y), .C(OR4_969_Y), .D(
        OR4_1159_Y), .Y(OR4_1761_Y));
    OR4 OR4_2834 (.A(\B_DOUT_TEMPR60[15] ), .B(\B_DOUT_TEMPR61[15] ), 
        .C(\B_DOUT_TEMPR62[15] ), .D(\B_DOUT_TEMPR63[15] ), .Y(
        OR4_2834_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%46%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R46C2 (
        .A_DOUT({nc24570, nc24571, nc24572, nc24573, nc24574, nc24575, 
        nc24576, nc24577, nc24578, nc24579, nc24580, nc24581, nc24582, 
        nc24583, nc24584, \A_DOUT_TEMPR46[14] , \A_DOUT_TEMPR46[13] , 
        \A_DOUT_TEMPR46[12] , \A_DOUT_TEMPR46[11] , 
        \A_DOUT_TEMPR46[10] }), .B_DOUT({nc24585, nc24586, nc24587, 
        nc24588, nc24589, nc24590, nc24591, nc24592, nc24593, nc24594, 
        nc24595, nc24596, nc24597, nc24598, nc24599, 
        \B_DOUT_TEMPR46[14] , \B_DOUT_TEMPR46[13] , 
        \B_DOUT_TEMPR46[12] , \B_DOUT_TEMPR46[11] , 
        \B_DOUT_TEMPR46[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[46][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%88%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R88C7 (
        .A_DOUT({nc24600, nc24601, nc24602, nc24603, nc24604, nc24605, 
        nc24606, nc24607, nc24608, nc24609, nc24610, nc24611, nc24612, 
        nc24613, nc24614, \A_DOUT_TEMPR88[39] , \A_DOUT_TEMPR88[38] , 
        \A_DOUT_TEMPR88[37] , \A_DOUT_TEMPR88[36] , 
        \A_DOUT_TEMPR88[35] }), .B_DOUT({nc24615, nc24616, nc24617, 
        nc24618, nc24619, nc24620, nc24621, nc24622, nc24623, nc24624, 
        nc24625, nc24626, nc24627, nc24628, nc24629, 
        \B_DOUT_TEMPR88[39] , \B_DOUT_TEMPR88[38] , 
        \B_DOUT_TEMPR88[37] , \B_DOUT_TEMPR88[36] , 
        \B_DOUT_TEMPR88[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[88][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1304 (.A(\A_DOUT_TEMPR95[27] ), .B(\A_DOUT_TEMPR96[27] ), 
        .C(\A_DOUT_TEMPR97[27] ), .D(\A_DOUT_TEMPR98[27] ), .Y(
        OR4_1304_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%40%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R40C6 (
        .A_DOUT({nc24630, nc24631, nc24632, nc24633, nc24634, nc24635, 
        nc24636, nc24637, nc24638, nc24639, nc24640, nc24641, nc24642, 
        nc24643, nc24644, \A_DOUT_TEMPR40[34] , \A_DOUT_TEMPR40[33] , 
        \A_DOUT_TEMPR40[32] , \A_DOUT_TEMPR40[31] , 
        \A_DOUT_TEMPR40[30] }), .B_DOUT({nc24645, nc24646, nc24647, 
        nc24648, nc24649, nc24650, nc24651, nc24652, nc24653, nc24654, 
        nc24655, nc24656, nc24657, nc24658, nc24659, 
        \B_DOUT_TEMPR40[34] , \B_DOUT_TEMPR40[33] , 
        \B_DOUT_TEMPR40[32] , \B_DOUT_TEMPR40[31] , 
        \B_DOUT_TEMPR40[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[40][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1244 (.A(\B_DOUT_TEMPR99[21] ), .B(\B_DOUT_TEMPR100[21] ), 
        .C(\B_DOUT_TEMPR101[21] ), .D(\B_DOUT_TEMPR102[21] ), .Y(
        OR4_1244_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%40%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R40C5 (
        .A_DOUT({nc24660, nc24661, nc24662, nc24663, nc24664, nc24665, 
        nc24666, nc24667, nc24668, nc24669, nc24670, nc24671, nc24672, 
        nc24673, nc24674, \A_DOUT_TEMPR40[29] , \A_DOUT_TEMPR40[28] , 
        \A_DOUT_TEMPR40[27] , \A_DOUT_TEMPR40[26] , 
        \A_DOUT_TEMPR40[25] }), .B_DOUT({nc24675, nc24676, nc24677, 
        nc24678, nc24679, nc24680, nc24681, nc24682, nc24683, nc24684, 
        nc24685, nc24686, nc24687, nc24688, nc24689, 
        \B_DOUT_TEMPR40[29] , \B_DOUT_TEMPR40[28] , 
        \B_DOUT_TEMPR40[27] , \B_DOUT_TEMPR40[26] , 
        \B_DOUT_TEMPR40[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[40][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2485 (.A(\B_DOUT_TEMPR36[0] ), .B(\B_DOUT_TEMPR37[0] ), .C(
        \B_DOUT_TEMPR38[0] ), .D(\B_DOUT_TEMPR39[0] ), .Y(OR4_2485_Y));
    OR4 OR4_2796 (.A(\B_DOUT_TEMPR111[16] ), .B(\B_DOUT_TEMPR112[16] ), 
        .C(\B_DOUT_TEMPR113[16] ), .D(\B_DOUT_TEMPR114[16] ), .Y(
        OR4_2796_Y));
    OR4 OR4_1834 (.A(\A_DOUT_TEMPR68[22] ), .B(\A_DOUT_TEMPR69[22] ), 
        .C(\A_DOUT_TEMPR70[22] ), .D(\A_DOUT_TEMPR71[22] ), .Y(
        OR4_1834_Y));
    OR4 OR4_2051 (.A(OR4_906_Y), .B(OR4_86_Y), .C(OR4_2575_Y), .D(
        OR4_2027_Y), .Y(OR4_2051_Y));
    OR2 OR2_35 (.A(\B_DOUT_TEMPR72[22] ), .B(\B_DOUT_TEMPR73[22] ), .Y(
        OR2_35_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[7]  (.A(CFG3_2_Y), .B(CFG3_16_Y)
        , .Y(\BLKY2[7] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%61%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R61C2 (
        .A_DOUT({nc24690, nc24691, nc24692, nc24693, nc24694, nc24695, 
        nc24696, nc24697, nc24698, nc24699, nc24700, nc24701, nc24702, 
        nc24703, nc24704, \A_DOUT_TEMPR61[14] , \A_DOUT_TEMPR61[13] , 
        \A_DOUT_TEMPR61[12] , \A_DOUT_TEMPR61[11] , 
        \A_DOUT_TEMPR61[10] }), .B_DOUT({nc24705, nc24706, nc24707, 
        nc24708, nc24709, nc24710, nc24711, nc24712, nc24713, nc24714, 
        nc24715, nc24716, nc24717, nc24718, nc24719, 
        \B_DOUT_TEMPR61[14] , \B_DOUT_TEMPR61[13] , 
        \B_DOUT_TEMPR61[12] , \B_DOUT_TEMPR61[11] , 
        \B_DOUT_TEMPR61[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[61][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_388 (.A(OR4_1979_Y), .B(OR4_81_Y), .C(OR4_444_Y), .D(
        OR4_753_Y), .Y(OR4_388_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%93%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R93C7 (
        .A_DOUT({nc24720, nc24721, nc24722, nc24723, nc24724, nc24725, 
        nc24726, nc24727, nc24728, nc24729, nc24730, nc24731, nc24732, 
        nc24733, nc24734, \A_DOUT_TEMPR93[39] , \A_DOUT_TEMPR93[38] , 
        \A_DOUT_TEMPR93[37] , \A_DOUT_TEMPR93[36] , 
        \A_DOUT_TEMPR93[35] }), .B_DOUT({nc24735, nc24736, nc24737, 
        nc24738, nc24739, nc24740, nc24741, nc24742, nc24743, nc24744, 
        nc24745, nc24746, nc24747, nc24748, nc24749, 
        \B_DOUT_TEMPR93[39] , \B_DOUT_TEMPR93[38] , 
        \B_DOUT_TEMPR93[37] , \B_DOUT_TEMPR93[36] , 
        \B_DOUT_TEMPR93[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[93][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_785 (.A(OR4_795_Y), .B(OR4_2769_Y), .C(OR4_333_Y), .D(
        OR4_2578_Y), .Y(OR4_785_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%13%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R13C1 (
        .A_DOUT({nc24750, nc24751, nc24752, nc24753, nc24754, nc24755, 
        nc24756, nc24757, nc24758, nc24759, nc24760, nc24761, nc24762, 
        nc24763, nc24764, \A_DOUT_TEMPR13[9] , \A_DOUT_TEMPR13[8] , 
        \A_DOUT_TEMPR13[7] , \A_DOUT_TEMPR13[6] , \A_DOUT_TEMPR13[5] })
        , .B_DOUT({nc24765, nc24766, nc24767, nc24768, nc24769, 
        nc24770, nc24771, nc24772, nc24773, nc24774, nc24775, nc24776, 
        nc24777, nc24778, nc24779, \B_DOUT_TEMPR13[9] , 
        \B_DOUT_TEMPR13[8] , \B_DOUT_TEMPR13[7] , \B_DOUT_TEMPR13[6] , 
        \B_DOUT_TEMPR13[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1043 (.A(\B_DOUT_TEMPR103[25] ), .B(\B_DOUT_TEMPR104[25] ), 
        .C(\B_DOUT_TEMPR105[25] ), .D(\B_DOUT_TEMPR106[25] ), .Y(
        OR4_1043_Y));
    OR4 \OR4_A_DOUT[16]  (.A(OR4_1541_Y), .B(OR4_2173_Y), .C(OR4_975_Y)
        , .D(OR4_989_Y), .Y(A_DOUT[16]));
    OR4 OR4_599 (.A(\B_DOUT_TEMPR103[39] ), .B(\B_DOUT_TEMPR104[39] ), 
        .C(\B_DOUT_TEMPR105[39] ), .D(\B_DOUT_TEMPR106[39] ), .Y(
        OR4_599_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENA[2]  (.A(A_WBYTE_EN[1]), .B(
        A_WEN), .Y(\WBYTEENA[2] ));
    OR4 OR4_1641 (.A(\A_DOUT_TEMPR91[20] ), .B(\A_DOUT_TEMPR92[20] ), 
        .C(\A_DOUT_TEMPR93[20] ), .D(\A_DOUT_TEMPR94[20] ), .Y(
        OR4_1641_Y));
    OR4 OR4_2740 (.A(OR4_538_Y), .B(OR4_953_Y), .C(OR4_1654_Y), .D(
        OR4_2475_Y), .Y(OR4_2740_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%4%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R4C7 (
        .A_DOUT({nc24780, nc24781, nc24782, nc24783, nc24784, nc24785, 
        nc24786, nc24787, nc24788, nc24789, nc24790, nc24791, nc24792, 
        nc24793, nc24794, \A_DOUT_TEMPR4[39] , \A_DOUT_TEMPR4[38] , 
        \A_DOUT_TEMPR4[37] , \A_DOUT_TEMPR4[36] , \A_DOUT_TEMPR4[35] })
        , .B_DOUT({nc24795, nc24796, nc24797, nc24798, nc24799, 
        nc24800, nc24801, nc24802, nc24803, nc24804, nc24805, nc24806, 
        nc24807, nc24808, nc24809, \B_DOUT_TEMPR4[39] , 
        \B_DOUT_TEMPR4[38] , \B_DOUT_TEMPR4[37] , \B_DOUT_TEMPR4[36] , 
        \B_DOUT_TEMPR4[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2786 (.A(OR4_1290_Y), .B(OR4_290_Y), .C(OR4_509_Y), .D(
        OR4_295_Y), .Y(OR4_2786_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%23%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R23C3 (
        .A_DOUT({nc24810, nc24811, nc24812, nc24813, nc24814, nc24815, 
        nc24816, nc24817, nc24818, nc24819, nc24820, nc24821, nc24822, 
        nc24823, nc24824, \A_DOUT_TEMPR23[19] , \A_DOUT_TEMPR23[18] , 
        \A_DOUT_TEMPR23[17] , \A_DOUT_TEMPR23[16] , 
        \A_DOUT_TEMPR23[15] }), .B_DOUT({nc24825, nc24826, nc24827, 
        nc24828, nc24829, nc24830, nc24831, nc24832, nc24833, nc24834, 
        nc24835, nc24836, nc24837, nc24838, nc24839, 
        \B_DOUT_TEMPR23[19] , \B_DOUT_TEMPR23[18] , 
        \B_DOUT_TEMPR23[17] , \B_DOUT_TEMPR23[16] , 
        \B_DOUT_TEMPR23[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1743 (.A(\B_DOUT_TEMPR0[9] ), .B(\B_DOUT_TEMPR1[9] ), .C(
        \B_DOUT_TEMPR2[9] ), .D(\B_DOUT_TEMPR3[9] ), .Y(OR4_1743_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%4%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R4C2 (
        .A_DOUT({nc24840, nc24841, nc24842, nc24843, nc24844, nc24845, 
        nc24846, nc24847, nc24848, nc24849, nc24850, nc24851, nc24852, 
        nc24853, nc24854, \A_DOUT_TEMPR4[14] , \A_DOUT_TEMPR4[13] , 
        \A_DOUT_TEMPR4[12] , \A_DOUT_TEMPR4[11] , \A_DOUT_TEMPR4[10] })
        , .B_DOUT({nc24855, nc24856, nc24857, nc24858, nc24859, 
        nc24860, nc24861, nc24862, nc24863, nc24864, nc24865, nc24866, 
        nc24867, nc24868, nc24869, \B_DOUT_TEMPR4[14] , 
        \B_DOUT_TEMPR4[13] , \B_DOUT_TEMPR4[12] , \B_DOUT_TEMPR4[11] , 
        \B_DOUT_TEMPR4[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[4][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1089 (.A(\B_DOUT_TEMPR75[1] ), .B(\B_DOUT_TEMPR76[1] ), .C(
        \B_DOUT_TEMPR77[1] ), .D(\B_DOUT_TEMPR78[1] ), .Y(OR4_1089_Y));
    OR4 OR4_453 (.A(\B_DOUT_TEMPR8[21] ), .B(\B_DOUT_TEMPR9[21] ), .C(
        \B_DOUT_TEMPR10[21] ), .D(\B_DOUT_TEMPR11[21] ), .Y(OR4_453_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_16 (.A(B_BLK_EN), .B(B_ADDR[18]), .C(
        B_ADDR[17]), .Y(CFG3_16_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%25%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R25C3 (
        .A_DOUT({nc24870, nc24871, nc24872, nc24873, nc24874, nc24875, 
        nc24876, nc24877, nc24878, nc24879, nc24880, nc24881, nc24882, 
        nc24883, nc24884, \A_DOUT_TEMPR25[19] , \A_DOUT_TEMPR25[18] , 
        \A_DOUT_TEMPR25[17] , \A_DOUT_TEMPR25[16] , 
        \A_DOUT_TEMPR25[15] }), .B_DOUT({nc24885, nc24886, nc24887, 
        nc24888, nc24889, nc24890, nc24891, nc24892, nc24893, nc24894, 
        nc24895, nc24896, nc24897, nc24898, nc24899, 
        \B_DOUT_TEMPR25[19] , \B_DOUT_TEMPR25[18] , 
        \B_DOUT_TEMPR25[17] , \B_DOUT_TEMPR25[16] , 
        \B_DOUT_TEMPR25[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[25][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1463 (.A(\B_DOUT_TEMPR44[26] ), .B(\B_DOUT_TEMPR45[26] ), 
        .C(\B_DOUT_TEMPR46[26] ), .D(\B_DOUT_TEMPR47[26] ), .Y(
        OR4_1463_Y));
    OR4 OR4_1145 (.A(\B_DOUT_TEMPR64[30] ), .B(\B_DOUT_TEMPR65[30] ), 
        .C(\B_DOUT_TEMPR66[30] ), .D(\B_DOUT_TEMPR67[30] ), .Y(
        OR4_1145_Y));
    OR4 OR4_2502 (.A(\A_DOUT_TEMPR99[13] ), .B(\A_DOUT_TEMPR100[13] ), 
        .C(\A_DOUT_TEMPR101[13] ), .D(\A_DOUT_TEMPR102[13] ), .Y(
        OR4_2502_Y));
    OR4 OR4_9 (.A(OR4_466_Y), .B(OR4_2704_Y), .C(OR4_1646_Y), .D(
        OR4_1962_Y), .Y(OR4_9_Y));
    OR4 OR4_1589 (.A(OR4_1588_Y), .B(OR4_1976_Y), .C(OR4_2748_Y), .D(
        OR4_506_Y), .Y(OR4_1589_Y));
    OR4 OR4_1475 (.A(\B_DOUT_TEMPR4[21] ), .B(\B_DOUT_TEMPR5[21] ), .C(
        \B_DOUT_TEMPR6[21] ), .D(\B_DOUT_TEMPR7[21] ), .Y(OR4_1475_Y));
    OR4 OR4_988 (.A(OR4_364_Y), .B(OR4_1679_Y), .C(OR4_1351_Y), .D(
        OR4_2373_Y), .Y(OR4_988_Y));
    OR4 OR4_86 (.A(OR4_162_Y), .B(OR4_1249_Y), .C(OR4_2958_Y), .D(
        OR4_1339_Y), .Y(OR4_86_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%109%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R109C0 (
        .A_DOUT({nc24900, nc24901, nc24902, nc24903, nc24904, nc24905, 
        nc24906, nc24907, nc24908, nc24909, nc24910, nc24911, nc24912, 
        nc24913, nc24914, \A_DOUT_TEMPR109[4] , \A_DOUT_TEMPR109[3] , 
        \A_DOUT_TEMPR109[2] , \A_DOUT_TEMPR109[1] , 
        \A_DOUT_TEMPR109[0] }), .B_DOUT({nc24915, nc24916, nc24917, 
        nc24918, nc24919, nc24920, nc24921, nc24922, nc24923, nc24924, 
        nc24925, nc24926, nc24927, nc24928, nc24929, 
        \B_DOUT_TEMPR109[4] , \B_DOUT_TEMPR109[3] , 
        \B_DOUT_TEMPR109[2] , \B_DOUT_TEMPR109[1] , 
        \B_DOUT_TEMPR109[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[109][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%81%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R81C1 (
        .A_DOUT({nc24930, nc24931, nc24932, nc24933, nc24934, nc24935, 
        nc24936, nc24937, nc24938, nc24939, nc24940, nc24941, nc24942, 
        nc24943, nc24944, \A_DOUT_TEMPR81[9] , \A_DOUT_TEMPR81[8] , 
        \A_DOUT_TEMPR81[7] , \A_DOUT_TEMPR81[6] , \A_DOUT_TEMPR81[5] })
        , .B_DOUT({nc24945, nc24946, nc24947, nc24948, nc24949, 
        nc24950, nc24951, nc24952, nc24953, nc24954, nc24955, nc24956, 
        nc24957, nc24958, nc24959, \B_DOUT_TEMPR81[9] , 
        \B_DOUT_TEMPR81[8] , \B_DOUT_TEMPR81[7] , \B_DOUT_TEMPR81[6] , 
        \B_DOUT_TEMPR81[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[81][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_470 (.A(\B_DOUT_TEMPR32[34] ), .B(\B_DOUT_TEMPR33[34] ), 
        .C(\B_DOUT_TEMPR34[34] ), .D(\B_DOUT_TEMPR35[34] ), .Y(
        OR4_470_Y));
    OR4 OR4_3028 (.A(\A_DOUT_TEMPR20[0] ), .B(\A_DOUT_TEMPR21[0] ), .C(
        \A_DOUT_TEMPR22[0] ), .D(\A_DOUT_TEMPR23[0] ), .Y(OR4_3028_Y));
    OR4 OR4_2014 (.A(OR4_3002_Y), .B(OR4_1187_Y), .C(OR4_1792_Y), .D(
        OR4_1011_Y), .Y(OR4_2014_Y));
    OR4 OR4_2016 (.A(\A_DOUT_TEMPR48[9] ), .B(\A_DOUT_TEMPR49[9] ), .C(
        \A_DOUT_TEMPR50[9] ), .D(\A_DOUT_TEMPR51[9] ), .Y(OR4_2016_Y));
    OR4 OR4_1129 (.A(\A_DOUT_TEMPR87[17] ), .B(\A_DOUT_TEMPR88[17] ), 
        .C(\A_DOUT_TEMPR89[17] ), .D(\A_DOUT_TEMPR90[17] ), .Y(
        OR4_1129_Y));
    OR4 OR4_1382 (.A(OR4_2221_Y), .B(OR4_2542_Y), .C(OR4_1124_Y), .D(
        OR4_2028_Y), .Y(OR4_1382_Y));
    OR4 OR4_1041 (.A(\A_DOUT_TEMPR103[17] ), .B(\A_DOUT_TEMPR104[17] ), 
        .C(\A_DOUT_TEMPR105[17] ), .D(\A_DOUT_TEMPR106[17] ), .Y(
        OR4_1041_Y));
    OR4 OR4_322 (.A(\B_DOUT_TEMPR60[19] ), .B(\B_DOUT_TEMPR61[19] ), 
        .C(\B_DOUT_TEMPR62[19] ), .D(\B_DOUT_TEMPR63[19] ), .Y(
        OR4_322_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%56%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R56C0 (
        .A_DOUT({nc24960, nc24961, nc24962, nc24963, nc24964, nc24965, 
        nc24966, nc24967, nc24968, nc24969, nc24970, nc24971, nc24972, 
        nc24973, nc24974, \A_DOUT_TEMPR56[4] , \A_DOUT_TEMPR56[3] , 
        \A_DOUT_TEMPR56[2] , \A_DOUT_TEMPR56[1] , \A_DOUT_TEMPR56[0] })
        , .B_DOUT({nc24975, nc24976, nc24977, nc24978, nc24979, 
        nc24980, nc24981, nc24982, nc24983, nc24984, nc24985, nc24986, 
        nc24987, nc24988, nc24989, \B_DOUT_TEMPR56[4] , 
        \B_DOUT_TEMPR56[3] , \B_DOUT_TEMPR56[2] , \B_DOUT_TEMPR56[1] , 
        \B_DOUT_TEMPR56[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[56][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2368 (.A(\B_DOUT_TEMPR52[20] ), .B(\B_DOUT_TEMPR53[20] ), 
        .C(\B_DOUT_TEMPR54[20] ), .D(\B_DOUT_TEMPR55[20] ), .Y(
        OR4_2368_Y));
    OR4 OR4_2347 (.A(\B_DOUT_TEMPR52[12] ), .B(\B_DOUT_TEMPR53[12] ), 
        .C(\B_DOUT_TEMPR54[12] ), .D(\B_DOUT_TEMPR55[12] ), .Y(
        OR4_2347_Y));
    OR4 OR4_188 (.A(\A_DOUT_TEMPR0[2] ), .B(\A_DOUT_TEMPR1[2] ), .C(
        \A_DOUT_TEMPR2[2] ), .D(\A_DOUT_TEMPR3[2] ), .Y(OR4_188_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%62%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R62C3 (
        .A_DOUT({nc24990, nc24991, nc24992, nc24993, nc24994, nc24995, 
        nc24996, nc24997, nc24998, nc24999, nc25000, nc25001, nc25002, 
        nc25003, nc25004, \A_DOUT_TEMPR62[19] , \A_DOUT_TEMPR62[18] , 
        \A_DOUT_TEMPR62[17] , \A_DOUT_TEMPR62[16] , 
        \A_DOUT_TEMPR62[15] }), .B_DOUT({nc25005, nc25006, nc25007, 
        nc25008, nc25009, nc25010, nc25011, nc25012, nc25013, nc25014, 
        nc25015, nc25016, nc25017, nc25018, nc25019, 
        \B_DOUT_TEMPR62[19] , \B_DOUT_TEMPR62[18] , 
        \B_DOUT_TEMPR62[17] , \B_DOUT_TEMPR62[16] , 
        \B_DOUT_TEMPR62[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[62][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2242 (.A(\B_DOUT_TEMPR48[0] ), .B(\B_DOUT_TEMPR49[0] ), .C(
        \B_DOUT_TEMPR50[0] ), .D(\B_DOUT_TEMPR51[0] ), .Y(OR4_2242_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%101%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R101C1 (
        .A_DOUT({nc25020, nc25021, nc25022, nc25023, nc25024, nc25025, 
        nc25026, nc25027, nc25028, nc25029, nc25030, nc25031, nc25032, 
        nc25033, nc25034, \A_DOUT_TEMPR101[9] , \A_DOUT_TEMPR101[8] , 
        \A_DOUT_TEMPR101[7] , \A_DOUT_TEMPR101[6] , 
        \A_DOUT_TEMPR101[5] }), .B_DOUT({nc25035, nc25036, nc25037, 
        nc25038, nc25039, nc25040, nc25041, nc25042, nc25043, nc25044, 
        nc25045, nc25046, nc25047, nc25048, nc25049, 
        \B_DOUT_TEMPR101[9] , \B_DOUT_TEMPR101[8] , 
        \B_DOUT_TEMPR101[7] , \B_DOUT_TEMPR101[6] , 
        \B_DOUT_TEMPR101[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[101][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1400 (.A(\A_DOUT_TEMPR87[21] ), .B(\A_DOUT_TEMPR88[21] ), 
        .C(\A_DOUT_TEMPR89[21] ), .D(\A_DOUT_TEMPR90[21] ), .Y(
        OR4_1400_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%48%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R48C5 (
        .A_DOUT({nc25050, nc25051, nc25052, nc25053, nc25054, nc25055, 
        nc25056, nc25057, nc25058, nc25059, nc25060, nc25061, nc25062, 
        nc25063, nc25064, \A_DOUT_TEMPR48[29] , \A_DOUT_TEMPR48[28] , 
        \A_DOUT_TEMPR48[27] , \A_DOUT_TEMPR48[26] , 
        \A_DOUT_TEMPR48[25] }), .B_DOUT({nc25065, nc25066, nc25067, 
        nc25068, nc25069, nc25070, nc25071, nc25072, nc25073, nc25074, 
        nc25075, nc25076, nc25077, nc25078, nc25079, 
        \B_DOUT_TEMPR48[29] , \B_DOUT_TEMPR48[28] , 
        \B_DOUT_TEMPR48[27] , \B_DOUT_TEMPR48[26] , 
        \B_DOUT_TEMPR48[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[48][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%60%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R60C3 (
        .A_DOUT({nc25080, nc25081, nc25082, nc25083, nc25084, nc25085, 
        nc25086, nc25087, nc25088, nc25089, nc25090, nc25091, nc25092, 
        nc25093, nc25094, \A_DOUT_TEMPR60[19] , \A_DOUT_TEMPR60[18] , 
        \A_DOUT_TEMPR60[17] , \A_DOUT_TEMPR60[16] , 
        \A_DOUT_TEMPR60[15] }), .B_DOUT({nc25095, nc25096, nc25097, 
        nc25098, nc25099, nc25100, nc25101, nc25102, nc25103, nc25104, 
        nc25105, nc25106, nc25107, nc25108, nc25109, 
        \B_DOUT_TEMPR60[19] , \B_DOUT_TEMPR60[18] , 
        \B_DOUT_TEMPR60[17] , \B_DOUT_TEMPR60[16] , 
        \B_DOUT_TEMPR60[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[60][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%93%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R93C0 (
        .A_DOUT({nc25110, nc25111, nc25112, nc25113, nc25114, nc25115, 
        nc25116, nc25117, nc25118, nc25119, nc25120, nc25121, nc25122, 
        nc25123, nc25124, \A_DOUT_TEMPR93[4] , \A_DOUT_TEMPR93[3] , 
        \A_DOUT_TEMPR93[2] , \A_DOUT_TEMPR93[1] , \A_DOUT_TEMPR93[0] })
        , .B_DOUT({nc25125, nc25126, nc25127, nc25128, nc25129, 
        nc25130, nc25131, nc25132, nc25133, nc25134, nc25135, nc25136, 
        nc25137, nc25138, nc25139, \B_DOUT_TEMPR93[4] , 
        \B_DOUT_TEMPR93[3] , \B_DOUT_TEMPR93[2] , \B_DOUT_TEMPR93[1] , 
        \B_DOUT_TEMPR93[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[93][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1776 (.A(OR4_2522_Y), .B(OR4_1179_Y), .C(OR4_597_Y), .D(
        OR4_1918_Y), .Y(OR4_1776_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%108%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R108C2 (
        .A_DOUT({nc25140, nc25141, nc25142, nc25143, nc25144, nc25145, 
        nc25146, nc25147, nc25148, nc25149, nc25150, nc25151, nc25152, 
        nc25153, nc25154, \A_DOUT_TEMPR108[14] , \A_DOUT_TEMPR108[13] , 
        \A_DOUT_TEMPR108[12] , \A_DOUT_TEMPR108[11] , 
        \A_DOUT_TEMPR108[10] }), .B_DOUT({nc25155, nc25156, nc25157, 
        nc25158, nc25159, nc25160, nc25161, nc25162, nc25163, nc25164, 
        nc25165, nc25166, nc25167, nc25168, nc25169, 
        \B_DOUT_TEMPR108[14] , \B_DOUT_TEMPR108[13] , 
        \B_DOUT_TEMPR108[12] , \B_DOUT_TEMPR108[11] , 
        \B_DOUT_TEMPR108[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[108][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%20%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R20C1 (
        .A_DOUT({nc25170, nc25171, nc25172, nc25173, nc25174, nc25175, 
        nc25176, nc25177, nc25178, nc25179, nc25180, nc25181, nc25182, 
        nc25183, nc25184, \A_DOUT_TEMPR20[9] , \A_DOUT_TEMPR20[8] , 
        \A_DOUT_TEMPR20[7] , \A_DOUT_TEMPR20[6] , \A_DOUT_TEMPR20[5] })
        , .B_DOUT({nc25185, nc25186, nc25187, nc25188, nc25189, 
        nc25190, nc25191, nc25192, nc25193, nc25194, nc25195, nc25196, 
        nc25197, nc25198, nc25199, \B_DOUT_TEMPR20[9] , 
        \B_DOUT_TEMPR20[8] , \B_DOUT_TEMPR20[7] , \B_DOUT_TEMPR20[6] , 
        \B_DOUT_TEMPR20[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_389 (.A(\B_DOUT_TEMPR16[21] ), .B(\B_DOUT_TEMPR17[21] ), 
        .C(\B_DOUT_TEMPR18[21] ), .D(\B_DOUT_TEMPR19[21] ), .Y(
        OR4_389_Y));
    OR4 OR4_2029 (.A(\B_DOUT_TEMPR0[25] ), .B(\B_DOUT_TEMPR1[25] ), .C(
        \B_DOUT_TEMPR2[25] ), .D(\B_DOUT_TEMPR3[25] ), .Y(OR4_2029_Y));
    OR2 OR2_21 (.A(\A_DOUT_TEMPR72[36] ), .B(\A_DOUT_TEMPR73[36] ), .Y(
        OR2_21_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%114%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R114C6 (
        .A_DOUT({nc25200, nc25201, nc25202, nc25203, nc25204, nc25205, 
        nc25206, nc25207, nc25208, nc25209, nc25210, nc25211, nc25212, 
        nc25213, nc25214, \A_DOUT_TEMPR114[34] , \A_DOUT_TEMPR114[33] , 
        \A_DOUT_TEMPR114[32] , \A_DOUT_TEMPR114[31] , 
        \A_DOUT_TEMPR114[30] }), .B_DOUT({nc25215, nc25216, nc25217, 
        nc25218, nc25219, nc25220, nc25221, nc25222, nc25223, nc25224, 
        nc25225, nc25226, nc25227, nc25228, nc25229, 
        \B_DOUT_TEMPR114[34] , \B_DOUT_TEMPR114[33] , 
        \B_DOUT_TEMPR114[32] , \B_DOUT_TEMPR114[31] , 
        \B_DOUT_TEMPR114[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[114][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2313 (.A(\A_DOUT_TEMPR44[13] ), .B(\A_DOUT_TEMPR45[13] ), 
        .C(\A_DOUT_TEMPR46[13] ), .D(\A_DOUT_TEMPR47[13] ), .Y(
        OR4_2313_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENB[6]  (.A(B_WBYTE_EN[3]), .B(
        B_WEN), .Y(\WBYTEENB[6] ));
    OR4 OR4_2529 (.A(\B_DOUT_TEMPR8[6] ), .B(\B_DOUT_TEMPR9[6] ), .C(
        \B_DOUT_TEMPR10[6] ), .D(\B_DOUT_TEMPR11[6] ), .Y(OR4_2529_Y));
    OR4 OR4_2597 (.A(\A_DOUT_TEMPR103[7] ), .B(\A_DOUT_TEMPR104[7] ), 
        .C(\A_DOUT_TEMPR105[7] ), .D(\A_DOUT_TEMPR106[7] ), .Y(
        OR4_2597_Y));
    OR4 OR4_1205 (.A(\A_DOUT_TEMPR16[33] ), .B(\A_DOUT_TEMPR17[33] ), 
        .C(\A_DOUT_TEMPR18[33] ), .D(\A_DOUT_TEMPR19[33] ), .Y(
        OR4_1205_Y));
    OR4 OR4_2335 (.A(OR4_768_Y), .B(OR4_1919_Y), .C(OR4_2263_Y), .D(
        OR4_2744_Y), .Y(OR4_2335_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%66%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R66C6 (
        .A_DOUT({nc25230, nc25231, nc25232, nc25233, nc25234, nc25235, 
        nc25236, nc25237, nc25238, nc25239, nc25240, nc25241, nc25242, 
        nc25243, nc25244, \A_DOUT_TEMPR66[34] , \A_DOUT_TEMPR66[33] , 
        \A_DOUT_TEMPR66[32] , \A_DOUT_TEMPR66[31] , 
        \A_DOUT_TEMPR66[30] }), .B_DOUT({nc25245, nc25246, nc25247, 
        nc25248, nc25249, nc25250, nc25251, nc25252, nc25253, nc25254, 
        nc25255, nc25256, nc25257, nc25258, nc25259, 
        \B_DOUT_TEMPR66[34] , \B_DOUT_TEMPR66[33] , 
        \B_DOUT_TEMPR66[32] , \B_DOUT_TEMPR66[31] , 
        \B_DOUT_TEMPR66[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[66][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1585 (.A(\A_DOUT_TEMPR44[18] ), .B(\A_DOUT_TEMPR45[18] ), 
        .C(\A_DOUT_TEMPR46[18] ), .D(\A_DOUT_TEMPR47[18] ), .Y(
        OR4_1585_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%41%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R41C7 (
        .A_DOUT({nc25260, nc25261, nc25262, nc25263, nc25264, nc25265, 
        nc25266, nc25267, nc25268, nc25269, nc25270, nc25271, nc25272, 
        nc25273, nc25274, \A_DOUT_TEMPR41[39] , \A_DOUT_TEMPR41[38] , 
        \A_DOUT_TEMPR41[37] , \A_DOUT_TEMPR41[36] , 
        \A_DOUT_TEMPR41[35] }), .B_DOUT({nc25275, nc25276, nc25277, 
        nc25278, nc25279, nc25280, nc25281, nc25282, nc25283, nc25284, 
        nc25285, nc25286, nc25287, nc25288, nc25289, 
        \B_DOUT_TEMPR41[39] , \B_DOUT_TEMPR41[38] , 
        \B_DOUT_TEMPR41[37] , \B_DOUT_TEMPR41[36] , 
        \B_DOUT_TEMPR41[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[41][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%97%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R97C7 (
        .A_DOUT({nc25290, nc25291, nc25292, nc25293, nc25294, nc25295, 
        nc25296, nc25297, nc25298, nc25299, nc25300, nc25301, nc25302, 
        nc25303, nc25304, \A_DOUT_TEMPR97[39] , \A_DOUT_TEMPR97[38] , 
        \A_DOUT_TEMPR97[37] , \A_DOUT_TEMPR97[36] , 
        \A_DOUT_TEMPR97[35] }), .B_DOUT({nc25305, nc25306, nc25307, 
        nc25308, nc25309, nc25310, nc25311, nc25312, nc25313, nc25314, 
        nc25315, nc25316, nc25317, nc25318, nc25319, 
        \B_DOUT_TEMPR97[39] , \B_DOUT_TEMPR97[38] , 
        \B_DOUT_TEMPR97[37] , \B_DOUT_TEMPR97[36] , 
        \B_DOUT_TEMPR97[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[97][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2444 (.A(\A_DOUT_TEMPR64[8] ), .B(\A_DOUT_TEMPR65[8] ), .C(
        \A_DOUT_TEMPR66[8] ), .D(\A_DOUT_TEMPR67[8] ), .Y(OR4_2444_Y));
    OR4 OR4_2000 (.A(\B_DOUT_TEMPR36[23] ), .B(\B_DOUT_TEMPR37[23] ), 
        .C(\B_DOUT_TEMPR38[23] ), .D(\B_DOUT_TEMPR39[23] ), .Y(
        OR4_2000_Y));
    OR4 OR4_3003 (.A(\B_DOUT_TEMPR52[1] ), .B(\B_DOUT_TEMPR53[1] ), .C(
        \B_DOUT_TEMPR54[1] ), .D(\B_DOUT_TEMPR55[1] ), .Y(OR4_3003_Y));
    OR4 OR4_525 (.A(\B_DOUT_TEMPR28[34] ), .B(\B_DOUT_TEMPR29[34] ), 
        .C(\B_DOUT_TEMPR30[34] ), .D(\B_DOUT_TEMPR31[34] ), .Y(
        OR4_525_Y));
    OR4 OR4_179 (.A(\B_DOUT_TEMPR24[8] ), .B(\B_DOUT_TEMPR25[8] ), .C(
        \B_DOUT_TEMPR26[8] ), .D(\B_DOUT_TEMPR27[8] ), .Y(OR4_179_Y));
    OR4 OR4_213 (.A(\B_DOUT_TEMPR95[8] ), .B(\B_DOUT_TEMPR96[8] ), .C(
        \B_DOUT_TEMPR97[8] ), .D(\B_DOUT_TEMPR98[8] ), .Y(OR4_213_Y));
    OR4 OR4_400 (.A(\A_DOUT_TEMPR103[30] ), .B(\A_DOUT_TEMPR104[30] ), 
        .C(\A_DOUT_TEMPR105[30] ), .D(\A_DOUT_TEMPR106[30] ), .Y(
        OR4_400_Y));
    OR4 OR4_1335 (.A(\B_DOUT_TEMPR68[18] ), .B(\B_DOUT_TEMPR69[18] ), 
        .C(\B_DOUT_TEMPR70[18] ), .D(\B_DOUT_TEMPR71[18] ), .Y(
        OR4_1335_Y));
    OR4 OR4_2322 (.A(\A_DOUT_TEMPR4[24] ), .B(\A_DOUT_TEMPR5[24] ), .C(
        \A_DOUT_TEMPR6[24] ), .D(\A_DOUT_TEMPR7[24] ), .Y(OR4_2322_Y));
    OR2 OR2_39 (.A(\A_DOUT_TEMPR72[21] ), .B(\A_DOUT_TEMPR73[21] ), .Y(
        OR2_39_Y));
    OR4 OR4_311 (.A(OR4_790_Y), .B(OR4_3032_Y), .C(OR4_1992_Y), .D(
        OR4_2280_Y), .Y(OR4_311_Y));
    OR4 OR4_815 (.A(\B_DOUT_TEMPR20[8] ), .B(\B_DOUT_TEMPR21[8] ), .C(
        \B_DOUT_TEMPR22[8] ), .D(\B_DOUT_TEMPR23[8] ), .Y(OR4_815_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%9%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R9C3 (
        .A_DOUT({nc25320, nc25321, nc25322, nc25323, nc25324, nc25325, 
        nc25326, nc25327, nc25328, nc25329, nc25330, nc25331, nc25332, 
        nc25333, nc25334, \A_DOUT_TEMPR9[19] , \A_DOUT_TEMPR9[18] , 
        \A_DOUT_TEMPR9[17] , \A_DOUT_TEMPR9[16] , \A_DOUT_TEMPR9[15] })
        , .B_DOUT({nc25335, nc25336, nc25337, nc25338, nc25339, 
        nc25340, nc25341, nc25342, nc25343, nc25344, nc25345, nc25346, 
        nc25347, nc25348, nc25349, \B_DOUT_TEMPR9[19] , 
        \B_DOUT_TEMPR9[18] , \B_DOUT_TEMPR9[17] , \B_DOUT_TEMPR9[16] , 
        \B_DOUT_TEMPR9[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_113 (.A(\A_DOUT_TEMPR32[34] ), .B(\A_DOUT_TEMPR33[34] ), 
        .C(\A_DOUT_TEMPR34[34] ), .D(\A_DOUT_TEMPR35[34] ), .Y(
        OR4_113_Y));
    OR4 OR4_282 (.A(\A_DOUT_TEMPR40[24] ), .B(\A_DOUT_TEMPR41[24] ), 
        .C(\A_DOUT_TEMPR42[24] ), .D(\A_DOUT_TEMPR43[24] ), .Y(
        OR4_282_Y));
    OR4 OR4_2971 (.A(\A_DOUT_TEMPR115[5] ), .B(\A_DOUT_TEMPR116[5] ), 
        .C(\A_DOUT_TEMPR117[5] ), .D(\A_DOUT_TEMPR118[5] ), .Y(
        OR4_2971_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%9%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R9C1 (
        .A_DOUT({nc25350, nc25351, nc25352, nc25353, nc25354, nc25355, 
        nc25356, nc25357, nc25358, nc25359, nc25360, nc25361, nc25362, 
        nc25363, nc25364, \A_DOUT_TEMPR9[9] , \A_DOUT_TEMPR9[8] , 
        \A_DOUT_TEMPR9[7] , \A_DOUT_TEMPR9[6] , \A_DOUT_TEMPR9[5] }), 
        .B_DOUT({nc25365, nc25366, nc25367, nc25368, nc25369, nc25370, 
        nc25371, nc25372, nc25373, nc25374, nc25375, nc25376, nc25377, 
        nc25378, nc25379, \B_DOUT_TEMPR9[9] , \B_DOUT_TEMPR9[8] , 
        \B_DOUT_TEMPR9[7] , \B_DOUT_TEMPR9[6] , \B_DOUT_TEMPR9[5] }), 
        .DB_DETECT(), .SB_CORRECT(), .ACCESS_BUSY(\ACCESS_BUSY[9][1] ), 
        .A_ADDR({A_ADDR[11], A_ADDR[10], A_ADDR[9], A_ADDR[8], 
        A_ADDR[7], A_ADDR[6], A_ADDR[5], A_ADDR[4], A_ADDR[3], 
        A_ADDR[2], A_ADDR[1], A_ADDR[0], GND, GND}), .A_BLK_EN({
        \BLKX2[2] , \BLKX1[0] , A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, A_DIN[9], A_DIN[8], A_DIN[7], A_DIN[6], 
        A_DIN[5]}), .A_REN(A_REN), .A_WEN({GND, \WBYTEENA[2] }), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({B_ADDR[11], B_ADDR[10], B_ADDR[9], B_ADDR[8], 
        B_ADDR[7], B_ADDR[6], B_ADDR[5], B_ADDR[4], B_ADDR[3], 
        B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, GND}), .B_BLK_EN({
        \BLKY2[2] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(B_CLK), .B_DIN({
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], B_DIN[6], 
        B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] }), 
        .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%0%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R0C3 (
        .A_DOUT({nc25380, nc25381, nc25382, nc25383, nc25384, nc25385, 
        nc25386, nc25387, nc25388, nc25389, nc25390, nc25391, nc25392, 
        nc25393, nc25394, \A_DOUT_TEMPR0[19] , \A_DOUT_TEMPR0[18] , 
        \A_DOUT_TEMPR0[17] , \A_DOUT_TEMPR0[16] , \A_DOUT_TEMPR0[15] })
        , .B_DOUT({nc25395, nc25396, nc25397, nc25398, nc25399, 
        nc25400, nc25401, nc25402, nc25403, nc25404, nc25405, nc25406, 
        nc25407, nc25408, nc25409, \B_DOUT_TEMPR0[19] , 
        \B_DOUT_TEMPR0[18] , \B_DOUT_TEMPR0[17] , \B_DOUT_TEMPR0[16] , 
        \B_DOUT_TEMPR0[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[0][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2587 (.A(\B_DOUT_TEMPR95[24] ), .B(\B_DOUT_TEMPR96[24] ), 
        .C(\B_DOUT_TEMPR97[24] ), .D(\B_DOUT_TEMPR98[24] ), .Y(
        OR4_2587_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%54%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R54C2 (
        .A_DOUT({nc25410, nc25411, nc25412, nc25413, nc25414, nc25415, 
        nc25416, nc25417, nc25418, nc25419, nc25420, nc25421, nc25422, 
        nc25423, nc25424, \A_DOUT_TEMPR54[14] , \A_DOUT_TEMPR54[13] , 
        \A_DOUT_TEMPR54[12] , \A_DOUT_TEMPR54[11] , 
        \A_DOUT_TEMPR54[10] }), .B_DOUT({nc25425, nc25426, nc25427, 
        nc25428, nc25429, nc25430, nc25431, nc25432, nc25433, nc25434, 
        nc25435, nc25436, nc25437, nc25438, nc25439, 
        \B_DOUT_TEMPR54[14] , \B_DOUT_TEMPR54[13] , 
        \B_DOUT_TEMPR54[12] , \B_DOUT_TEMPR54[11] , 
        \B_DOUT_TEMPR54[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[54][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2465 (.A(OR4_471_Y), .B(OR4_1642_Y), .C(OR4_2727_Y), .D(
        OR4_526_Y), .Y(OR4_2465_Y));
    OR4 \OR4_B_DOUT[24]  (.A(OR4_1469_Y), .B(OR4_501_Y), .C(OR4_348_Y), 
        .D(OR4_125_Y), .Y(B_DOUT[24]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%11%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R11C2 (
        .A_DOUT({nc25440, nc25441, nc25442, nc25443, nc25444, nc25445, 
        nc25446, nc25447, nc25448, nc25449, nc25450, nc25451, nc25452, 
        nc25453, nc25454, \A_DOUT_TEMPR11[14] , \A_DOUT_TEMPR11[13] , 
        \A_DOUT_TEMPR11[12] , \A_DOUT_TEMPR11[11] , 
        \A_DOUT_TEMPR11[10] }), .B_DOUT({nc25455, nc25456, nc25457, 
        nc25458, nc25459, nc25460, nc25461, nc25462, nc25463, nc25464, 
        nc25465, nc25466, nc25467, nc25468, nc25469, 
        \B_DOUT_TEMPR11[14] , \B_DOUT_TEMPR11[13] , 
        \B_DOUT_TEMPR11[12] , \B_DOUT_TEMPR11[11] , 
        \B_DOUT_TEMPR11[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[11][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_342 (.A(\B_DOUT_TEMPR87[31] ), .B(\B_DOUT_TEMPR88[31] ), 
        .C(\B_DOUT_TEMPR89[31] ), .D(\B_DOUT_TEMPR90[31] ), .Y(
        OR4_342_Y));
    OR4 OR4_837 (.A(\B_DOUT_TEMPR52[38] ), .B(\B_DOUT_TEMPR53[38] ), 
        .C(\B_DOUT_TEMPR54[38] ), .D(\B_DOUT_TEMPR55[38] ), .Y(
        OR4_837_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%36%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R36C0 (
        .A_DOUT({nc25470, nc25471, nc25472, nc25473, nc25474, nc25475, 
        nc25476, nc25477, nc25478, nc25479, nc25480, nc25481, nc25482, 
        nc25483, nc25484, \A_DOUT_TEMPR36[4] , \A_DOUT_TEMPR36[3] , 
        \A_DOUT_TEMPR36[2] , \A_DOUT_TEMPR36[1] , \A_DOUT_TEMPR36[0] })
        , .B_DOUT({nc25485, nc25486, nc25487, nc25488, nc25489, 
        nc25490, nc25491, nc25492, nc25493, nc25494, nc25495, nc25496, 
        nc25497, nc25498, nc25499, \B_DOUT_TEMPR36[4] , 
        \B_DOUT_TEMPR36[3] , \B_DOUT_TEMPR36[2] , \B_DOUT_TEMPR36[1] , 
        \B_DOUT_TEMPR36[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1266 (.A(\A_DOUT_TEMPR75[37] ), .B(\A_DOUT_TEMPR76[37] ), 
        .C(\A_DOUT_TEMPR77[37] ), .D(\A_DOUT_TEMPR78[37] ), .Y(
        OR4_1266_Y));
    OR4 OR4_493 (.A(OR4_1634_Y), .B(OR4_2864_Y), .C(OR4_856_Y), .D(
        OR4_626_Y), .Y(OR4_493_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[6]  (.A(CFG3_19_Y), .B(
        CFG3_16_Y), .Y(\BLKY2[6] ));
    OR4 OR4_1988 (.A(\A_DOUT_TEMPR36[20] ), .B(\A_DOUT_TEMPR37[20] ), 
        .C(\A_DOUT_TEMPR38[20] ), .D(\A_DOUT_TEMPR39[20] ), .Y(
        OR4_1988_Y));
    OR4 OR4_1951 (.A(\A_DOUT_TEMPR28[26] ), .B(\A_DOUT_TEMPR29[26] ), 
        .C(\A_DOUT_TEMPR30[26] ), .D(\A_DOUT_TEMPR31[26] ), .Y(
        OR4_1951_Y));
    OR4 OR4_2525 (.A(OR4_823_Y), .B(OR4_2489_Y), .C(OR4_1936_Y), .D(
        OR4_205_Y), .Y(OR4_2525_Y));
    OR4 OR4_3001 (.A(\A_DOUT_TEMPR75[2] ), .B(\A_DOUT_TEMPR76[2] ), .C(
        \A_DOUT_TEMPR77[2] ), .D(\A_DOUT_TEMPR78[2] ), .Y(OR4_3001_Y));
    OR4 OR4_1822 (.A(OR4_2851_Y), .B(OR4_2017_Y), .C(OR4_1012_Y), .D(
        OR4_1303_Y), .Y(OR4_1822_Y));
    OR4 OR4_1615 (.A(\A_DOUT_TEMPR75[14] ), .B(\A_DOUT_TEMPR76[14] ), 
        .C(\A_DOUT_TEMPR77[14] ), .D(\A_DOUT_TEMPR78[14] ), .Y(
        OR4_1615_Y));
    OR4 OR4_712 (.A(\B_DOUT_TEMPR48[37] ), .B(\B_DOUT_TEMPR49[37] ), 
        .C(\B_DOUT_TEMPR50[37] ), .D(\B_DOUT_TEMPR51[37] ), .Y(
        OR4_712_Y));
    OR4 OR4_2406 (.A(OR4_2042_Y), .B(OR4_312_Y), .C(OR4_3023_Y), .D(
        OR4_1048_Y), .Y(OR4_2406_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%53%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R53C7 (
        .A_DOUT({nc25500, nc25501, nc25502, nc25503, nc25504, nc25505, 
        nc25506, nc25507, nc25508, nc25509, nc25510, nc25511, nc25512, 
        nc25513, nc25514, \A_DOUT_TEMPR53[39] , \A_DOUT_TEMPR53[38] , 
        \A_DOUT_TEMPR53[37] , \A_DOUT_TEMPR53[36] , 
        \A_DOUT_TEMPR53[35] }), .B_DOUT({nc25515, nc25516, nc25517, 
        nc25518, nc25519, nc25520, nc25521, nc25522, nc25523, nc25524, 
        nc25525, nc25526, nc25527, nc25528, nc25529, 
        \B_DOUT_TEMPR53[39] , \B_DOUT_TEMPR53[38] , 
        \B_DOUT_TEMPR53[37] , \B_DOUT_TEMPR53[36] , 
        \B_DOUT_TEMPR53[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[53][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_316 (.A(\A_DOUT_TEMPR75[32] ), .B(\A_DOUT_TEMPR76[32] ), 
        .C(\A_DOUT_TEMPR77[32] ), .D(\A_DOUT_TEMPR78[32] ), .Y(
        OR4_316_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%76%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R76C1 (
        .A_DOUT({nc25530, nc25531, nc25532, nc25533, nc25534, nc25535, 
        nc25536, nc25537, nc25538, nc25539, nc25540, nc25541, nc25542, 
        nc25543, nc25544, \A_DOUT_TEMPR76[9] , \A_DOUT_TEMPR76[8] , 
        \A_DOUT_TEMPR76[7] , \A_DOUT_TEMPR76[6] , \A_DOUT_TEMPR76[5] })
        , .B_DOUT({nc25545, nc25546, nc25547, nc25548, nc25549, 
        nc25550, nc25551, nc25552, nc25553, nc25554, nc25555, nc25556, 
        nc25557, nc25558, nc25559, \B_DOUT_TEMPR76[9] , 
        \B_DOUT_TEMPR76[8] , \B_DOUT_TEMPR76[7] , \B_DOUT_TEMPR76[6] , 
        \B_DOUT_TEMPR76[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[76][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2273 (.A(\A_DOUT_TEMPR60[30] ), .B(\A_DOUT_TEMPR61[30] ), 
        .C(\A_DOUT_TEMPR62[30] ), .D(\A_DOUT_TEMPR63[30] ), .Y(
        OR4_2273_Y));
    OR4 OR4_109 (.A(\A_DOUT_TEMPR52[3] ), .B(\A_DOUT_TEMPR53[3] ), .C(
        \A_DOUT_TEMPR54[3] ), .D(\A_DOUT_TEMPR55[3] ), .Y(OR4_109_Y));
    OR4 OR4_2766 (.A(\B_DOUT_TEMPR79[21] ), .B(\B_DOUT_TEMPR80[21] ), 
        .C(\B_DOUT_TEMPR81[21] ), .D(\B_DOUT_TEMPR82[21] ), .Y(
        OR4_2766_Y));
    OR4 OR4_7 (.A(OR4_1661_Y), .B(OR4_1961_Y), .C(OR4_1431_Y), .D(
        OR4_2526_Y), .Y(OR4_7_Y));
    OR4 OR4_771 (.A(OR4_1685_Y), .B(OR4_898_Y), .C(OR4_2924_Y), .D(
        OR4_146_Y), .Y(OR4_771_Y));
    OR4 OR4_2298 (.A(\A_DOUT_TEMPR20[29] ), .B(\A_DOUT_TEMPR21[29] ), 
        .C(\A_DOUT_TEMPR22[29] ), .D(\A_DOUT_TEMPR23[29] ), .Y(
        OR4_2298_Y));
    OR4 OR4_2244 (.A(OR4_2887_Y), .B(OR4_1494_Y), .C(OR4_968_Y), .D(
        OR4_2238_Y), .Y(OR4_2244_Y));
    OR4 OR4_1577 (.A(\A_DOUT_TEMPR20[36] ), .B(\A_DOUT_TEMPR21[36] ), 
        .C(\A_DOUT_TEMPR22[36] ), .D(\A_DOUT_TEMPR23[36] ), .Y(
        OR4_1577_Y));
    OR4 OR4_517 (.A(\B_DOUT_TEMPR103[1] ), .B(\B_DOUT_TEMPR104[1] ), 
        .C(\B_DOUT_TEMPR105[1] ), .D(\B_DOUT_TEMPR106[1] ), .Y(
        OR4_517_Y));
    OR4 OR4_545 (.A(\B_DOUT_TEMPR91[37] ), .B(\B_DOUT_TEMPR92[37] ), 
        .C(\B_DOUT_TEMPR93[37] ), .D(\B_DOUT_TEMPR94[37] ), .Y(
        OR4_545_Y));
    OR4 OR4_2705 (.A(\B_DOUT_TEMPR87[10] ), .B(\B_DOUT_TEMPR88[10] ), 
        .C(\B_DOUT_TEMPR89[10] ), .D(\B_DOUT_TEMPR90[10] ), .Y(
        OR4_2705_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%76%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R76C2 (
        .A_DOUT({nc25560, nc25561, nc25562, nc25563, nc25564, nc25565, 
        nc25566, nc25567, nc25568, nc25569, nc25570, nc25571, nc25572, 
        nc25573, nc25574, \A_DOUT_TEMPR76[14] , \A_DOUT_TEMPR76[13] , 
        \A_DOUT_TEMPR76[12] , \A_DOUT_TEMPR76[11] , 
        \A_DOUT_TEMPR76[10] }), .B_DOUT({nc25575, nc25576, nc25577, 
        nc25578, nc25579, nc25580, nc25581, nc25582, nc25583, nc25584, 
        nc25585, nc25586, nc25587, nc25588, nc25589, 
        \B_DOUT_TEMPR76[14] , \B_DOUT_TEMPR76[13] , 
        \B_DOUT_TEMPR76[12] , \B_DOUT_TEMPR76[11] , 
        \B_DOUT_TEMPR76[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[76][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1617 (.A(\B_DOUT_TEMPR83[28] ), .B(\B_DOUT_TEMPR84[28] ), 
        .C(\B_DOUT_TEMPR85[28] ), .D(\B_DOUT_TEMPR86[28] ), .Y(
        OR4_1617_Y));
    OR4 OR4_1606 (.A(\B_DOUT_TEMPR32[36] ), .B(\B_DOUT_TEMPR33[36] ), 
        .C(\B_DOUT_TEMPR34[36] ), .D(\B_DOUT_TEMPR35[36] ), .Y(
        OR4_1606_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%20%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R20C7 (
        .A_DOUT({nc25590, nc25591, nc25592, nc25593, nc25594, nc25595, 
        nc25596, nc25597, nc25598, nc25599, nc25600, nc25601, nc25602, 
        nc25603, nc25604, \A_DOUT_TEMPR20[39] , \A_DOUT_TEMPR20[38] , 
        \A_DOUT_TEMPR20[37] , \A_DOUT_TEMPR20[36] , 
        \A_DOUT_TEMPR20[35] }), .B_DOUT({nc25605, nc25606, nc25607, 
        nc25608, nc25609, nc25610, nc25611, nc25612, nc25613, nc25614, 
        nc25615, nc25616, nc25617, nc25618, nc25619, 
        \B_DOUT_TEMPR20[39] , \B_DOUT_TEMPR20[38] , 
        \B_DOUT_TEMPR20[37] , \B_DOUT_TEMPR20[36] , 
        \B_DOUT_TEMPR20[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%47%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R47C0 (
        .A_DOUT({nc25620, nc25621, nc25622, nc25623, nc25624, nc25625, 
        nc25626, nc25627, nc25628, nc25629, nc25630, nc25631, nc25632, 
        nc25633, nc25634, \A_DOUT_TEMPR47[4] , \A_DOUT_TEMPR47[3] , 
        \A_DOUT_TEMPR47[2] , \A_DOUT_TEMPR47[1] , \A_DOUT_TEMPR47[0] })
        , .B_DOUT({nc25635, nc25636, nc25637, nc25638, nc25639, 
        nc25640, nc25641, nc25642, nc25643, nc25644, nc25645, nc25646, 
        nc25647, nc25648, nc25649, \B_DOUT_TEMPR47[4] , 
        \B_DOUT_TEMPR47[3] , \B_DOUT_TEMPR47[2] , \B_DOUT_TEMPR47[1] , 
        \B_DOUT_TEMPR47[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%70%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R70C6 (
        .A_DOUT({nc25650, nc25651, nc25652, nc25653, nc25654, nc25655, 
        nc25656, nc25657, nc25658, nc25659, nc25660, nc25661, nc25662, 
        nc25663, nc25664, \A_DOUT_TEMPR70[34] , \A_DOUT_TEMPR70[33] , 
        \A_DOUT_TEMPR70[32] , \A_DOUT_TEMPR70[31] , 
        \A_DOUT_TEMPR70[30] }), .B_DOUT({nc25665, nc25666, nc25667, 
        nc25668, nc25669, nc25670, nc25671, nc25672, nc25673, nc25674, 
        nc25675, nc25676, nc25677, nc25678, nc25679, 
        \B_DOUT_TEMPR70[34] , \B_DOUT_TEMPR70[33] , 
        \B_DOUT_TEMPR70[32] , \B_DOUT_TEMPR70[31] , 
        \B_DOUT_TEMPR70[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[70][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_67 (.A(\B_DOUT_TEMPR72[33] ), .B(\B_DOUT_TEMPR73[33] ), .Y(
        OR2_67_Y));
    OR4 OR4_1100 (.A(\A_DOUT_TEMPR52[20] ), .B(\A_DOUT_TEMPR53[20] ), 
        .C(\A_DOUT_TEMPR54[20] ), .D(\A_DOUT_TEMPR55[20] ), .Y(
        OR4_1100_Y));
    OR4 OR4_1253 (.A(\B_DOUT_TEMPR91[36] ), .B(\B_DOUT_TEMPR92[36] ), 
        .C(\B_DOUT_TEMPR93[36] ), .D(\B_DOUT_TEMPR94[36] ), .Y(
        OR4_1253_Y));
    OR4 OR4_1623 (.A(\A_DOUT_TEMPR20[24] ), .B(\A_DOUT_TEMPR21[24] ), 
        .C(\A_DOUT_TEMPR22[24] ), .D(\A_DOUT_TEMPR23[24] ), .Y(
        OR4_1623_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%70%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R70C5 (
        .A_DOUT({nc25680, nc25681, nc25682, nc25683, nc25684, nc25685, 
        nc25686, nc25687, nc25688, nc25689, nc25690, nc25691, nc25692, 
        nc25693, nc25694, \A_DOUT_TEMPR70[29] , \A_DOUT_TEMPR70[28] , 
        \A_DOUT_TEMPR70[27] , \A_DOUT_TEMPR70[26] , 
        \A_DOUT_TEMPR70[25] }), .B_DOUT({nc25695, nc25696, nc25697, 
        nc25698, nc25699, nc25700, nc25701, nc25702, nc25703, nc25704, 
        nc25705, nc25706, nc25707, nc25708, nc25709, 
        \B_DOUT_TEMPR70[29] , \B_DOUT_TEMPR70[28] , 
        \B_DOUT_TEMPR70[27] , \B_DOUT_TEMPR70[26] , 
        \B_DOUT_TEMPR70[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[70][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2655 (.A(OR4_1968_Y), .B(OR4_2810_Y), .C(OR4_1840_Y), .D(
        OR4_1651_Y), .Y(OR4_2655_Y));
    OR4 OR4_2043 (.A(\B_DOUT_TEMPR64[25] ), .B(\B_DOUT_TEMPR65[25] ), 
        .C(\B_DOUT_TEMPR66[25] ), .D(\B_DOUT_TEMPR67[25] ), .Y(
        OR4_2043_Y));
    OR4 OR4_1187 (.A(\A_DOUT_TEMPR36[22] ), .B(\A_DOUT_TEMPR37[22] ), 
        .C(\A_DOUT_TEMPR38[22] ), .D(\A_DOUT_TEMPR39[22] ), .Y(
        OR4_1187_Y));
    OR4 OR4_1866 (.A(OR4_2053_Y), .B(OR4_1255_Y), .C(OR4_200_Y), .D(
        OR4_518_Y), .Y(OR4_1866_Y));
    OR4 OR4_2928 (.A(OR4_565_Y), .B(OR4_1746_Y), .C(OR4_2822_Y), .D(
        OR4_2405_Y), .Y(OR4_2928_Y));
    OR4 OR4_1929 (.A(\A_DOUT_TEMPR16[29] ), .B(\A_DOUT_TEMPR17[29] ), 
        .C(\A_DOUT_TEMPR18[29] ), .D(\A_DOUT_TEMPR19[29] ), .Y(
        OR4_1929_Y));
    OR4 OR4_1684 (.A(\A_DOUT_TEMPR91[21] ), .B(\A_DOUT_TEMPR92[21] ), 
        .C(\A_DOUT_TEMPR93[21] ), .D(\A_DOUT_TEMPR94[21] ), .Y(
        OR4_1684_Y));
    OR4 OR4_872 (.A(\A_DOUT_TEMPR4[8] ), .B(\A_DOUT_TEMPR5[8] ), .C(
        \A_DOUT_TEMPR6[8] ), .D(\A_DOUT_TEMPR7[8] ), .Y(OR4_872_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%34%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R34C2 (
        .A_DOUT({nc25710, nc25711, nc25712, nc25713, nc25714, nc25715, 
        nc25716, nc25717, nc25718, nc25719, nc25720, nc25721, nc25722, 
        nc25723, nc25724, \A_DOUT_TEMPR34[14] , \A_DOUT_TEMPR34[13] , 
        \A_DOUT_TEMPR34[12] , \A_DOUT_TEMPR34[11] , 
        \A_DOUT_TEMPR34[10] }), .B_DOUT({nc25725, nc25726, nc25727, 
        nc25728, nc25729, nc25730, nc25731, nc25732, nc25733, nc25734, 
        nc25735, nc25736, nc25737, nc25738, nc25739, 
        \B_DOUT_TEMPR34[14] , \B_DOUT_TEMPR34[13] , 
        \B_DOUT_TEMPR34[12] , \B_DOUT_TEMPR34[11] , 
        \B_DOUT_TEMPR34[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[34][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2288 (.A(\B_DOUT_TEMPR103[14] ), .B(\B_DOUT_TEMPR104[14] ), 
        .C(\B_DOUT_TEMPR105[14] ), .D(\B_DOUT_TEMPR106[14] ), .Y(
        OR4_2288_Y));
    OR2 OR2_17 (.A(\A_DOUT_TEMPR72[0] ), .B(\A_DOUT_TEMPR73[0] ), .Y(
        OR2_17_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%12%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R12C3 (
        .A_DOUT({nc25740, nc25741, nc25742, nc25743, nc25744, nc25745, 
        nc25746, nc25747, nc25748, nc25749, nc25750, nc25751, nc25752, 
        nc25753, nc25754, \A_DOUT_TEMPR12[19] , \A_DOUT_TEMPR12[18] , 
        \A_DOUT_TEMPR12[17] , \A_DOUT_TEMPR12[16] , 
        \A_DOUT_TEMPR12[15] }), .B_DOUT({nc25755, nc25756, nc25757, 
        nc25758, nc25759, nc25760, nc25761, nc25762, nc25763, nc25764, 
        nc25765, nc25766, nc25767, nc25768, nc25769, 
        \B_DOUT_TEMPR12[19] , \B_DOUT_TEMPR12[18] , 
        \B_DOUT_TEMPR12[17] , \B_DOUT_TEMPR12[16] , 
        \B_DOUT_TEMPR12[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[12][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2641 (.A(\A_DOUT_TEMPR75[13] ), .B(\A_DOUT_TEMPR76[13] ), 
        .C(\A_DOUT_TEMPR77[13] ), .D(\A_DOUT_TEMPR78[13] ), .Y(
        OR4_2641_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%10%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R10C3 (
        .A_DOUT({nc25770, nc25771, nc25772, nc25773, nc25774, nc25775, 
        nc25776, nc25777, nc25778, nc25779, nc25780, nc25781, nc25782, 
        nc25783, nc25784, \A_DOUT_TEMPR10[19] , \A_DOUT_TEMPR10[18] , 
        \A_DOUT_TEMPR10[17] , \A_DOUT_TEMPR10[16] , 
        \A_DOUT_TEMPR10[15] }), .B_DOUT({nc25785, nc25786, nc25787, 
        nc25788, nc25789, nc25790, nc25791, nc25792, nc25793, nc25794, 
        nc25795, nc25796, nc25797, nc25798, nc25799, 
        \B_DOUT_TEMPR10[19] , \B_DOUT_TEMPR10[18] , 
        \B_DOUT_TEMPR10[17] , \B_DOUT_TEMPR10[16] , 
        \B_DOUT_TEMPR10[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[10][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_450 (.A(\B_DOUT_TEMPR8[3] ), .B(\B_DOUT_TEMPR9[3] ), .C(
        \B_DOUT_TEMPR10[3] ), .D(\B_DOUT_TEMPR11[3] ), .Y(OR4_450_Y));
    OR4 OR4_2743 (.A(OR4_1883_Y), .B(OR4_1675_Y), .C(OR4_2552_Y), .D(
        OR4_708_Y), .Y(OR4_2743_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENA[6]  (.A(A_WBYTE_EN[3]), .B(
        A_WEN), .Y(\WBYTEENA[6] ));
    OR2 OR2_26 (.A(\B_DOUT_TEMPR72[30] ), .B(\B_DOUT_TEMPR73[30] ), .Y(
        OR2_26_Y));
    OR4 OR4_2145 (.A(OR4_436_Y), .B(OR4_728_Y), .C(OR4_2329_Y), .D(
        OR4_214_Y), .Y(OR4_2145_Y));
    OR4 OR4_701 (.A(OR4_2596_Y), .B(OR4_1598_Y), .C(OR4_1805_Y), .D(
        OR4_1609_Y), .Y(OR4_701_Y));
    OR4 OR4_2657 (.A(\A_DOUT_TEMPR107[35] ), .B(\A_DOUT_TEMPR108[35] ), 
        .C(\A_DOUT_TEMPR109[35] ), .D(\A_DOUT_TEMPR110[35] ), .Y(
        OR4_2657_Y));
    OR4 OR4_431 (.A(\B_DOUT_TEMPR12[14] ), .B(\B_DOUT_TEMPR13[14] ), 
        .C(\B_DOUT_TEMPR14[14] ), .D(\B_DOUT_TEMPR15[14] ), .Y(
        OR4_431_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%117%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R117C5 (
        .A_DOUT({nc25800, nc25801, nc25802, nc25803, nc25804, nc25805, 
        nc25806, nc25807, nc25808, nc25809, nc25810, nc25811, nc25812, 
        nc25813, nc25814, \A_DOUT_TEMPR117[29] , \A_DOUT_TEMPR117[28] , 
        \A_DOUT_TEMPR117[27] , \A_DOUT_TEMPR117[26] , 
        \A_DOUT_TEMPR117[25] }), .B_DOUT({nc25815, nc25816, nc25817, 
        nc25818, nc25819, nc25820, nc25821, nc25822, nc25823, nc25824, 
        nc25825, nc25826, nc25827, nc25828, nc25829, 
        \B_DOUT_TEMPR117[29] , \B_DOUT_TEMPR117[28] , 
        \B_DOUT_TEMPR117[27] , \B_DOUT_TEMPR117[26] , 
        \B_DOUT_TEMPR117[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[117][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%33%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R33C7 (
        .A_DOUT({nc25830, nc25831, nc25832, nc25833, nc25834, nc25835, 
        nc25836, nc25837, nc25838, nc25839, nc25840, nc25841, nc25842, 
        nc25843, nc25844, \A_DOUT_TEMPR33[39] , \A_DOUT_TEMPR33[38] , 
        \A_DOUT_TEMPR33[37] , \A_DOUT_TEMPR33[36] , 
        \A_DOUT_TEMPR33[35] }), .B_DOUT({nc25845, nc25846, nc25847, 
        nc25848, nc25849, nc25850, nc25851, nc25852, nc25853, nc25854, 
        nc25855, nc25856, nc25857, nc25858, nc25859, 
        \B_DOUT_TEMPR33[39] , \B_DOUT_TEMPR33[38] , 
        \B_DOUT_TEMPR33[37] , \B_DOUT_TEMPR33[36] , 
        \B_DOUT_TEMPR33[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[33][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1724 (.A(\B_DOUT_TEMPR56[21] ), .B(\B_DOUT_TEMPR57[21] ), 
        .C(\B_DOUT_TEMPR58[21] ), .D(\B_DOUT_TEMPR59[21] ), .Y(
        OR4_1724_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%16%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R16C6 (
        .A_DOUT({nc25860, nc25861, nc25862, nc25863, nc25864, nc25865, 
        nc25866, nc25867, nc25868, nc25869, nc25870, nc25871, nc25872, 
        nc25873, nc25874, \A_DOUT_TEMPR16[34] , \A_DOUT_TEMPR16[33] , 
        \A_DOUT_TEMPR16[32] , \A_DOUT_TEMPR16[31] , 
        \A_DOUT_TEMPR16[30] }), .B_DOUT({nc25875, nc25876, nc25877, 
        nc25878, nc25879, nc25880, nc25881, nc25882, nc25883, nc25884, 
        nc25885, nc25886, nc25887, nc25888, nc25889, 
        \B_DOUT_TEMPR16[34] , \B_DOUT_TEMPR16[33] , 
        \B_DOUT_TEMPR16[32] , \B_DOUT_TEMPR16[31] , 
        \B_DOUT_TEMPR16[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%53%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R53C0 (
        .A_DOUT({nc25890, nc25891, nc25892, nc25893, nc25894, nc25895, 
        nc25896, nc25897, nc25898, nc25899, nc25900, nc25901, nc25902, 
        nc25903, nc25904, \A_DOUT_TEMPR53[4] , \A_DOUT_TEMPR53[3] , 
        \A_DOUT_TEMPR53[2] , \A_DOUT_TEMPR53[1] , \A_DOUT_TEMPR53[0] })
        , .B_DOUT({nc25905, nc25906, nc25907, nc25908, nc25909, 
        nc25910, nc25911, nc25912, nc25913, nc25914, nc25915, nc25916, 
        nc25917, nc25918, nc25919, \B_DOUT_TEMPR53[4] , 
        \B_DOUT_TEMPR53[3] , \B_DOUT_TEMPR53[2] , \B_DOUT_TEMPR53[1] , 
        \B_DOUT_TEMPR53[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[53][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[13] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1421 (.A(OR4_2283_Y), .B(OR4_1475_Y), .C(OR4_453_Y), .D(
        OR4_752_Y), .Y(OR4_1421_Y));
    OR4 OR4_263 (.A(\A_DOUT_TEMPR107[16] ), .B(\A_DOUT_TEMPR108[16] ), 
        .C(\A_DOUT_TEMPR109[16] ), .D(\A_DOUT_TEMPR110[16] ), .Y(
        OR4_263_Y));
    OR4 OR4_2041 (.A(\A_DOUT_TEMPR20[18] ), .B(\A_DOUT_TEMPR21[18] ), 
        .C(\A_DOUT_TEMPR22[18] ), .D(\A_DOUT_TEMPR23[18] ), .Y(
        OR4_2041_Y));
    OR4 OR4_1760 (.A(\B_DOUT_TEMPR8[28] ), .B(\B_DOUT_TEMPR9[28] ), .C(
        \B_DOUT_TEMPR10[28] ), .D(\B_DOUT_TEMPR11[28] ), .Y(OR4_1760_Y)
        );
    OR4 OR4_2127 (.A(\B_DOUT_TEMPR12[38] ), .B(\B_DOUT_TEMPR13[38] ), 
        .C(\B_DOUT_TEMPR14[38] ), .D(\B_DOUT_TEMPR15[38] ), .Y(
        OR4_2127_Y));
    OR4 OR4_361 (.A(\A_DOUT_TEMPR111[26] ), .B(\A_DOUT_TEMPR112[26] ), 
        .C(\A_DOUT_TEMPR113[26] ), .D(\A_DOUT_TEMPR114[26] ), .Y(
        OR4_361_Y));
    OR2 OR2_60 (.A(\B_DOUT_TEMPR72[12] ), .B(\B_DOUT_TEMPR73[12] ), .Y(
        OR2_60_Y));
    OR4 OR4_1278 (.A(OR4_1929_Y), .B(OR4_2298_Y), .C(OR4_32_Y), .D(
        OR4_836_Y), .Y(OR4_1278_Y));
    OR4 OR4_2624 (.A(\B_DOUT_TEMPR28[18] ), .B(\B_DOUT_TEMPR29[18] ), 
        .C(\B_DOUT_TEMPR30[18] ), .D(\B_DOUT_TEMPR31[18] ), .Y(
        OR4_2624_Y));
    OR4 OR4_865 (.A(\A_DOUT_TEMPR0[22] ), .B(\A_DOUT_TEMPR1[22] ), .C(
        \A_DOUT_TEMPR2[22] ), .D(\A_DOUT_TEMPR3[22] ), .Y(OR4_865_Y));
    OR4 OR4_163 (.A(OR4_1056_Y), .B(OR4_850_Y), .C(OR4_1697_Y), .D(
        OR4_2930_Y), .Y(OR4_163_Y));
    OR4 OR4_802 (.A(\B_DOUT_TEMPR36[5] ), .B(\B_DOUT_TEMPR37[5] ), .C(
        \B_DOUT_TEMPR38[5] ), .D(\B_DOUT_TEMPR39[5] ), .Y(OR4_802_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%57%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R57C7 (
        .A_DOUT({nc25920, nc25921, nc25922, nc25923, nc25924, nc25925, 
        nc25926, nc25927, nc25928, nc25929, nc25930, nc25931, nc25932, 
        nc25933, nc25934, \A_DOUT_TEMPR57[39] , \A_DOUT_TEMPR57[38] , 
        \A_DOUT_TEMPR57[37] , \A_DOUT_TEMPR57[36] , 
        \A_DOUT_TEMPR57[35] }), .B_DOUT({nc25935, nc25936, nc25937, 
        nc25938, nc25939, nc25940, nc25941, nc25942, nc25943, nc25944, 
        nc25945, nc25946, nc25947, nc25948, nc25949, 
        \B_DOUT_TEMPR57[39] , \B_DOUT_TEMPR57[38] , 
        \B_DOUT_TEMPR57[37] , \B_DOUT_TEMPR57[36] , 
        \B_DOUT_TEMPR57[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[57][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_328 (.A(\B_DOUT_TEMPR36[36] ), .B(\B_DOUT_TEMPR37[36] ), 
        .C(\B_DOUT_TEMPR38[36] ), .D(\B_DOUT_TEMPR39[36] ), .Y(
        OR4_328_Y));
    OR2 OR2_10 (.A(\B_DOUT_TEMPR72[39] ), .B(\B_DOUT_TEMPR73[39] ), .Y(
        OR2_10_Y));
    OR4 OR4_1314 (.A(\A_DOUT_TEMPR103[1] ), .B(\A_DOUT_TEMPR104[1] ), 
        .C(\A_DOUT_TEMPR105[1] ), .D(\A_DOUT_TEMPR106[1] ), .Y(
        OR4_1314_Y));
    OR4 OR4_1645 (.A(\B_DOUT_TEMPR115[38] ), .B(\B_DOUT_TEMPR116[38] ), 
        .C(\B_DOUT_TEMPR117[38] ), .D(\B_DOUT_TEMPR118[38] ), .Y(
        OR4_1645_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%106%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R106C1 (
        .A_DOUT({nc25950, nc25951, nc25952, nc25953, nc25954, nc25955, 
        nc25956, nc25957, nc25958, nc25959, nc25960, nc25961, nc25962, 
        nc25963, nc25964, \A_DOUT_TEMPR106[9] , \A_DOUT_TEMPR106[8] , 
        \A_DOUT_TEMPR106[7] , \A_DOUT_TEMPR106[6] , 
        \A_DOUT_TEMPR106[5] }), .B_DOUT({nc25965, nc25966, nc25967, 
        nc25968, nc25969, nc25970, nc25971, nc25972, nc25973, nc25974, 
        nc25975, nc25976, nc25977, nc25978, nc25979, 
        \B_DOUT_TEMPR106[9] , \B_DOUT_TEMPR106[8] , 
        \B_DOUT_TEMPR106[7] , \B_DOUT_TEMPR106[6] , 
        \B_DOUT_TEMPR106[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[106][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%118%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R118C5 (
        .A_DOUT({nc25980, nc25981, nc25982, nc25983, nc25984, nc25985, 
        nc25986, nc25987, nc25988, nc25989, nc25990, nc25991, nc25992, 
        nc25993, nc25994, \A_DOUT_TEMPR118[29] , \A_DOUT_TEMPR118[28] , 
        \A_DOUT_TEMPR118[27] , \A_DOUT_TEMPR118[26] , 
        \A_DOUT_TEMPR118[25] }), .B_DOUT({nc25995, nc25996, nc25997, 
        nc25998, nc25999, nc26000, nc26001, nc26002, nc26003, nc26004, 
        nc26005, nc26006, nc26007, nc26008, nc26009, 
        \B_DOUT_TEMPR118[29] , \B_DOUT_TEMPR118[28] , 
        \B_DOUT_TEMPR118[27] , \B_DOUT_TEMPR118[26] , 
        \B_DOUT_TEMPR118[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[118][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%83%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R83C2 (
        .A_DOUT({nc26010, nc26011, nc26012, nc26013, nc26014, nc26015, 
        nc26016, nc26017, nc26018, nc26019, nc26020, nc26021, nc26022, 
        nc26023, nc26024, \A_DOUT_TEMPR83[14] , \A_DOUT_TEMPR83[13] , 
        \A_DOUT_TEMPR83[12] , \A_DOUT_TEMPR83[11] , 
        \A_DOUT_TEMPR83[10] }), .B_DOUT({nc26025, nc26026, nc26027, 
        nc26028, nc26029, nc26030, nc26031, nc26032, nc26033, nc26034, 
        nc26035, nc26036, nc26037, nc26038, nc26039, 
        \B_DOUT_TEMPR83[14] , \B_DOUT_TEMPR83[13] , 
        \B_DOUT_TEMPR83[12] , \B_DOUT_TEMPR83[11] , 
        \B_DOUT_TEMPR83[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[83][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_725 (.A(\B_DOUT_TEMPR48[15] ), .B(\B_DOUT_TEMPR49[15] ), 
        .C(\B_DOUT_TEMPR50[15] ), .D(\B_DOUT_TEMPR51[15] ), .Y(
        OR4_725_Y));
    OR4 OR4_159 (.A(OR4_2943_Y), .B(OR4_799_Y), .C(OR4_445_Y), .D(
        OR4_1949_Y), .Y(OR4_159_Y));
    OR4 OR4_2567 (.A(\B_DOUT_TEMPR60[0] ), .B(\B_DOUT_TEMPR61[0] ), .C(
        \B_DOUT_TEMPR62[0] ), .D(\B_DOUT_TEMPR63[0] ), .Y(OR4_2567_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%66%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R66C0 (
        .A_DOUT({nc26040, nc26041, nc26042, nc26043, nc26044, nc26045, 
        nc26046, nc26047, nc26048, nc26049, nc26050, nc26051, nc26052, 
        nc26053, nc26054, \A_DOUT_TEMPR66[4] , \A_DOUT_TEMPR66[3] , 
        \A_DOUT_TEMPR66[2] , \A_DOUT_TEMPR66[1] , \A_DOUT_TEMPR66[0] })
        , .B_DOUT({nc26055, nc26056, nc26057, nc26058, nc26059, 
        nc26060, nc26061, nc26062, nc26063, nc26064, nc26065, nc26066, 
        nc26067, nc26068, nc26069, \B_DOUT_TEMPR66[4] , 
        \B_DOUT_TEMPR66[3] , \B_DOUT_TEMPR66[2] , \B_DOUT_TEMPR66[1] , 
        \B_DOUT_TEMPR66[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[66][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%22%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R22C0 (
        .A_DOUT({nc26070, nc26071, nc26072, nc26073, nc26074, nc26075, 
        nc26076, nc26077, nc26078, nc26079, nc26080, nc26081, nc26082, 
        nc26083, nc26084, \A_DOUT_TEMPR22[4] , \A_DOUT_TEMPR22[3] , 
        \A_DOUT_TEMPR22[2] , \A_DOUT_TEMPR22[1] , \A_DOUT_TEMPR22[0] })
        , .B_DOUT({nc26085, nc26086, nc26087, nc26088, nc26089, 
        nc26090, nc26091, nc26092, nc26093, nc26094, nc26095, nc26096, 
        nc26097, nc26098, nc26099, \B_DOUT_TEMPR22[4] , 
        \B_DOUT_TEMPR22[3] , \B_DOUT_TEMPR22[2] , \B_DOUT_TEMPR22[1] , 
        \B_DOUT_TEMPR22[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_716 (.A(\A_DOUT_TEMPR68[36] ), .B(\A_DOUT_TEMPR69[36] ), 
        .C(\A_DOUT_TEMPR70[36] ), .D(\A_DOUT_TEMPR71[36] ), .Y(
        OR4_716_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[1]  (.A(CFG3_8_Y), .B(CFG3_16_Y)
        , .Y(\BLKY2[1] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%78%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R78C5 (
        .A_DOUT({nc26100, nc26101, nc26102, nc26103, nc26104, nc26105, 
        nc26106, nc26107, nc26108, nc26109, nc26110, nc26111, nc26112, 
        nc26113, nc26114, \A_DOUT_TEMPR78[29] , \A_DOUT_TEMPR78[28] , 
        \A_DOUT_TEMPR78[27] , \A_DOUT_TEMPR78[26] , 
        \A_DOUT_TEMPR78[25] }), .B_DOUT({nc26115, nc26116, nc26117, 
        nc26118, nc26119, nc26120, nc26121, nc26122, nc26123, nc26124, 
        nc26125, nc26126, nc26127, nc26128, nc26129, 
        \B_DOUT_TEMPR78[29] , \B_DOUT_TEMPR78[28] , 
        \B_DOUT_TEMPR78[27] , \B_DOUT_TEMPR78[26] , 
        \B_DOUT_TEMPR78[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[78][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1924 (.A(\A_DOUT_TEMPR44[12] ), .B(\A_DOUT_TEMPR45[12] ), 
        .C(\A_DOUT_TEMPR46[12] ), .D(\A_DOUT_TEMPR47[12] ), .Y(
        OR4_1924_Y));
    OR4 OR4_1903 (.A(\A_DOUT_TEMPR16[1] ), .B(\A_DOUT_TEMPR17[1] ), .C(
        \A_DOUT_TEMPR18[1] ), .D(\A_DOUT_TEMPR19[1] ), .Y(OR4_1903_Y));
    OR4 OR4_2533 (.A(\B_DOUT_TEMPR60[9] ), .B(\B_DOUT_TEMPR61[9] ), .C(
        \B_DOUT_TEMPR62[9] ), .D(\B_DOUT_TEMPR63[9] ), .Y(OR4_2533_Y));
    OR4 OR4_2506 (.A(OR4_1517_Y), .B(OR4_1815_Y), .C(OR4_1447_Y), .D(
        OR4_1835_Y), .Y(OR4_2506_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%21%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R21C6 (
        .A_DOUT({nc26130, nc26131, nc26132, nc26133, nc26134, nc26135, 
        nc26136, nc26137, nc26138, nc26139, nc26140, nc26141, nc26142, 
        nc26143, nc26144, \A_DOUT_TEMPR21[34] , \A_DOUT_TEMPR21[33] , 
        \A_DOUT_TEMPR21[32] , \A_DOUT_TEMPR21[31] , 
        \A_DOUT_TEMPR21[30] }), .B_DOUT({nc26145, nc26146, nc26147, 
        nc26148, nc26149, nc26150, nc26151, nc26152, nc26153, nc26154, 
        nc26155, nc26156, nc26157, nc26158, nc26159, 
        \B_DOUT_TEMPR21[34] , \B_DOUT_TEMPR21[33] , 
        \B_DOUT_TEMPR21[32] , \B_DOUT_TEMPR21[31] , 
        \B_DOUT_TEMPR21[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1367 (.A(\A_DOUT_TEMPR87[20] ), .B(\A_DOUT_TEMPR88[20] ), 
        .C(\A_DOUT_TEMPR89[20] ), .D(\A_DOUT_TEMPR90[20] ), .Y(
        OR4_1367_Y));
    OR4 OR4_762 (.A(OR4_2781_Y), .B(OR4_1768_Y), .C(OR4_1981_Y), .D(
        OR4_1779_Y), .Y(OR4_762_Y));
    OR4 OR4_1262 (.A(\A_DOUT_TEMPR16[24] ), .B(\A_DOUT_TEMPR17[24] ), 
        .C(\A_DOUT_TEMPR18[24] ), .D(\A_DOUT_TEMPR19[24] ), .Y(
        OR4_1262_Y));
    OR4 OR4_1926 (.A(OR4_1189_Y), .B(OR4_1882_Y), .C(OR4_2583_Y), .D(
        OR4_2896_Y), .Y(OR4_1926_Y));
    OR4 OR4_1647 (.A(\B_DOUT_TEMPR103[28] ), .B(\B_DOUT_TEMPR104[28] ), 
        .C(\B_DOUT_TEMPR105[28] ), .D(\B_DOUT_TEMPR106[28] ), .Y(
        OR4_1647_Y));
    OR4 OR4_2707 (.A(\B_DOUT_TEMPR107[22] ), .B(\B_DOUT_TEMPR108[22] ), 
        .C(\B_DOUT_TEMPR109[22] ), .D(\B_DOUT_TEMPR110[22] ), .Y(
        OR4_2707_Y));
    OR4 OR4_777 (.A(\A_DOUT_TEMPR36[16] ), .B(\A_DOUT_TEMPR37[16] ), 
        .C(\A_DOUT_TEMPR38[16] ), .D(\A_DOUT_TEMPR39[16] ), .Y(
        OR4_777_Y));
    OR4 OR4_366 (.A(\A_DOUT_TEMPR12[26] ), .B(\A_DOUT_TEMPR13[26] ), 
        .C(\A_DOUT_TEMPR14[26] ), .D(\A_DOUT_TEMPR15[26] ), .Y(
        OR4_366_Y));
    OR4 OR4_2354 (.A(\A_DOUT_TEMPR103[14] ), .B(\A_DOUT_TEMPR104[14] ), 
        .C(\A_DOUT_TEMPR105[14] ), .D(\A_DOUT_TEMPR106[14] ), .Y(
        OR4_2354_Y));
    OR4 OR4_1533 (.A(\B_DOUT_TEMPR16[22] ), .B(\B_DOUT_TEMPR17[22] ), 
        .C(\B_DOUT_TEMPR18[22] ), .D(\B_DOUT_TEMPR19[22] ), .Y(
        OR4_1533_Y));
    OR4 OR4_2501 (.A(OR4_2479_Y), .B(OR4_1134_Y), .C(OR4_496_Y), .D(
        OR4_2874_Y), .Y(OR4_2501_Y));
    OR4 OR4_2133 (.A(\B_DOUT_TEMPR83[17] ), .B(\B_DOUT_TEMPR84[17] ), 
        .C(\B_DOUT_TEMPR85[17] ), .D(\B_DOUT_TEMPR86[17] ), .Y(
        OR4_2133_Y));
    OR4 OR4_373 (.A(OR4_2346_Y), .B(OR4_2661_Y), .C(OR4_1240_Y), .D(
        OR4_2127_Y), .Y(OR4_373_Y));
    OR4 OR4_928 (.A(\A_DOUT_TEMPR60[17] ), .B(\A_DOUT_TEMPR61[17] ), 
        .C(\A_DOUT_TEMPR62[17] ), .D(\A_DOUT_TEMPR63[17] ), .Y(
        OR4_928_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[3]  (.A(CFG3_20_Y), .B(
        CFG3_16_Y), .Y(\BLKY2[3] ));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%33%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R33C0 (
        .A_DOUT({nc26160, nc26161, nc26162, nc26163, nc26164, nc26165, 
        nc26166, nc26167, nc26168, nc26169, nc26170, nc26171, nc26172, 
        nc26173, nc26174, \A_DOUT_TEMPR33[4] , \A_DOUT_TEMPR33[3] , 
        \A_DOUT_TEMPR33[2] , \A_DOUT_TEMPR33[1] , \A_DOUT_TEMPR33[0] })
        , .B_DOUT({nc26175, nc26176, nc26177, nc26178, nc26179, 
        nc26180, nc26181, nc26182, nc26183, nc26184, nc26185, nc26186, 
        nc26187, nc26188, nc26189, \B_DOUT_TEMPR33[4] , 
        \B_DOUT_TEMPR33[3] , \B_DOUT_TEMPR33[2] , \B_DOUT_TEMPR33[1] , 
        \B_DOUT_TEMPR33[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[33][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[8] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%7%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R7C7 (
        .A_DOUT({nc26190, nc26191, nc26192, nc26193, nc26194, nc26195, 
        nc26196, nc26197, nc26198, nc26199, nc26200, nc26201, nc26202, 
        nc26203, nc26204, \A_DOUT_TEMPR7[39] , \A_DOUT_TEMPR7[38] , 
        \A_DOUT_TEMPR7[37] , \A_DOUT_TEMPR7[36] , \A_DOUT_TEMPR7[35] })
        , .B_DOUT({nc26205, nc26206, nc26207, nc26208, nc26209, 
        nc26210, nc26211, nc26212, nc26213, nc26214, nc26215, nc26216, 
        nc26217, nc26218, nc26219, \B_DOUT_TEMPR7[39] , 
        \B_DOUT_TEMPR7[38] , \B_DOUT_TEMPR7[37] , \B_DOUT_TEMPR7[36] , 
        \B_DOUT_TEMPR7[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[7][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2118 (.A(\B_DOUT_TEMPR16[3] ), .B(\B_DOUT_TEMPR17[3] ), .C(
        \B_DOUT_TEMPR18[3] ), .D(\B_DOUT_TEMPR19[3] ), .Y(OR4_2118_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%71%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R71C7 (
        .A_DOUT({nc26220, nc26221, nc26222, nc26223, nc26224, nc26225, 
        nc26226, nc26227, nc26228, nc26229, nc26230, nc26231, nc26232, 
        nc26233, nc26234, \A_DOUT_TEMPR71[39] , \A_DOUT_TEMPR71[38] , 
        \A_DOUT_TEMPR71[37] , \A_DOUT_TEMPR71[36] , 
        \A_DOUT_TEMPR71[35] }), .B_DOUT({nc26235, nc26236, nc26237, 
        nc26238, nc26239, nc26240, nc26241, nc26242, nc26243, nc26244, 
        nc26245, nc26246, nc26247, nc26248, nc26249, 
        \B_DOUT_TEMPR71[39] , \B_DOUT_TEMPR71[38] , 
        \B_DOUT_TEMPR71[37] , \B_DOUT_TEMPR71[36] , 
        \B_DOUT_TEMPR71[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[71][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%110%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R110C0 (
        .A_DOUT({nc26250, nc26251, nc26252, nc26253, nc26254, nc26255, 
        nc26256, nc26257, nc26258, nc26259, nc26260, nc26261, nc26262, 
        nc26263, nc26264, \A_DOUT_TEMPR110[4] , \A_DOUT_TEMPR110[3] , 
        \A_DOUT_TEMPR110[2] , \A_DOUT_TEMPR110[1] , 
        \A_DOUT_TEMPR110[0] }), .B_DOUT({nc26265, nc26266, nc26267, 
        nc26268, nc26269, nc26270, nc26271, nc26272, nc26273, nc26274, 
        nc26275, nc26276, nc26277, nc26278, nc26279, 
        \B_DOUT_TEMPR110[4] , \B_DOUT_TEMPR110[3] , 
        \B_DOUT_TEMPR110[2] , \B_DOUT_TEMPR110[1] , 
        \B_DOUT_TEMPR110[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[110][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_778 (.A(\B_DOUT_TEMPR16[7] ), .B(\B_DOUT_TEMPR17[7] ), .C(
        \B_DOUT_TEMPR18[7] ), .D(\B_DOUT_TEMPR19[7] ), .Y(OR4_778_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%89%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R89C4 (
        .A_DOUT({nc26280, nc26281, nc26282, nc26283, nc26284, nc26285, 
        nc26286, nc26287, nc26288, nc26289, nc26290, nc26291, nc26292, 
        nc26293, nc26294, \A_DOUT_TEMPR89[24] , \A_DOUT_TEMPR89[23] , 
        \A_DOUT_TEMPR89[22] , \A_DOUT_TEMPR89[21] , 
        \A_DOUT_TEMPR89[20] }), .B_DOUT({nc26295, nc26296, nc26297, 
        nc26298, nc26299, nc26300, nc26301, nc26302, nc26303, nc26304, 
        nc26305, nc26306, nc26307, nc26308, nc26309, 
        \B_DOUT_TEMPR89[24] , \B_DOUT_TEMPR89[23] , 
        \B_DOUT_TEMPR89[22] , \B_DOUT_TEMPR89[21] , 
        \B_DOUT_TEMPR89[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[89][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1680 (.A(\B_DOUT_TEMPR103[34] ), .B(\B_DOUT_TEMPR104[34] ), 
        .C(\B_DOUT_TEMPR105[34] ), .D(\B_DOUT_TEMPR106[34] ), .Y(
        OR4_1680_Y));
    OR4 OR4_1133 (.A(\B_DOUT_TEMPR60[23] ), .B(\B_DOUT_TEMPR61[23] ), 
        .C(\B_DOUT_TEMPR62[23] ), .D(\B_DOUT_TEMPR63[23] ), .Y(
        OR4_1133_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%49%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R49C6 (
        .A_DOUT({nc26310, nc26311, nc26312, nc26313, nc26314, nc26315, 
        nc26316, nc26317, nc26318, nc26319, nc26320, nc26321, nc26322, 
        nc26323, nc26324, \A_DOUT_TEMPR49[34] , \A_DOUT_TEMPR49[33] , 
        \A_DOUT_TEMPR49[32] , \A_DOUT_TEMPR49[31] , 
        \A_DOUT_TEMPR49[30] }), .B_DOUT({nc26325, nc26326, nc26327, 
        nc26328, nc26329, nc26330, nc26331, nc26332, nc26333, nc26334, 
        nc26335, nc26336, nc26337, nc26338, nc26339, 
        \B_DOUT_TEMPR49[34] , \B_DOUT_TEMPR49[33] , 
        \B_DOUT_TEMPR49[32] , \B_DOUT_TEMPR49[31] , 
        \B_DOUT_TEMPR49[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[49][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2032 (.A(\B_DOUT_TEMPR111[37] ), .B(\B_DOUT_TEMPR112[37] ), 
        .C(\B_DOUT_TEMPR113[37] ), .D(\B_DOUT_TEMPR114[37] ), .Y(
        OR4_2032_Y));
    OR4 OR4_1301 (.A(\A_DOUT_TEMPR95[20] ), .B(\A_DOUT_TEMPR96[20] ), 
        .C(\A_DOUT_TEMPR97[20] ), .D(\A_DOUT_TEMPR98[20] ), .Y(
        OR4_1301_Y));
    OR4 OR4_511 (.A(OR4_1425_Y), .B(OR4_182_Y), .C(OR4_2881_Y), .D(
        OR4_1289_Y), .Y(OR4_511_Y));
    OR4 OR4_673 (.A(\A_DOUT_TEMPR87[23] ), .B(\A_DOUT_TEMPR88[23] ), 
        .C(\A_DOUT_TEMPR89[23] ), .D(\A_DOUT_TEMPR90[23] ), .Y(
        OR4_673_Y));
    OR4 OR4_567 (.A(\B_DOUT_TEMPR0[1] ), .B(\B_DOUT_TEMPR1[1] ), .C(
        \B_DOUT_TEMPR2[1] ), .D(\B_DOUT_TEMPR3[1] ), .Y(OR4_567_Y));
    OR4 OR4_518 (.A(\A_DOUT_TEMPR12[28] ), .B(\A_DOUT_TEMPR13[28] ), 
        .C(\A_DOUT_TEMPR14[28] ), .D(\A_DOUT_TEMPR15[28] ), .Y(
        OR4_518_Y));
    OR4 OR4_3012 (.A(OR4_1106_Y), .B(OR4_2985_Y), .C(OR4_2543_Y), .D(
        OR4_1198_Y), .Y(OR4_3012_Y));
    OR4 OR4_1801 (.A(\A_DOUT_TEMPR44[20] ), .B(\A_DOUT_TEMPR45[20] ), 
        .C(\A_DOUT_TEMPR46[20] ), .D(\A_DOUT_TEMPR47[20] ), .Y(
        OR4_1801_Y));
    OR4 OR4_1088 (.A(\B_DOUT_TEMPR115[29] ), .B(\B_DOUT_TEMPR116[29] ), 
        .C(\B_DOUT_TEMPR117[29] ), .D(\B_DOUT_TEMPR118[29] ), .Y(
        OR4_1088_Y));
    OR4 OR4_1032 (.A(\B_DOUT_TEMPR68[1] ), .B(\B_DOUT_TEMPR69[1] ), .C(
        \B_DOUT_TEMPR70[1] ), .D(\B_DOUT_TEMPR71[1] ), .Y(OR4_1032_Y));
    OR4 \OR4_A_DOUT[14]  (.A(OR4_1782_Y), .B(OR4_396_Y), .C(OR4_580_Y), 
        .D(OR4_1817_Y), .Y(A_DOUT[14]));
    OR4 OR4_1464 (.A(\B_DOUT_TEMPR20[27] ), .B(\B_DOUT_TEMPR21[27] ), 
        .C(\B_DOUT_TEMPR22[27] ), .D(\B_DOUT_TEMPR23[27] ), .Y(
        OR4_1464_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%116%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R116C6 (
        .A_DOUT({nc26340, nc26341, nc26342, nc26343, nc26344, nc26345, 
        nc26346, nc26347, nc26348, nc26349, nc26350, nc26351, nc26352, 
        nc26353, nc26354, \A_DOUT_TEMPR116[34] , \A_DOUT_TEMPR116[33] , 
        \A_DOUT_TEMPR116[32] , \A_DOUT_TEMPR116[31] , 
        \A_DOUT_TEMPR116[30] }), .B_DOUT({nc26355, nc26356, nc26357, 
        nc26358, nc26359, nc26360, nc26361, nc26362, nc26363, nc26364, 
        nc26365, nc26366, nc26367, nc26368, nc26369, 
        \B_DOUT_TEMPR116[34] , \B_DOUT_TEMPR116[33] , 
        \B_DOUT_TEMPR116[32] , \B_DOUT_TEMPR116[31] , 
        \B_DOUT_TEMPR116[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[116][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[29] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[29] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_490 (.A(OR4_1262_Y), .B(OR4_1623_Y), .C(OR4_2362_Y), .D(
        OR4_138_Y), .Y(OR4_490_Y));
    OR4 OR4_128 (.A(\A_DOUT_TEMPR91[17] ), .B(\A_DOUT_TEMPR92[17] ), 
        .C(\A_DOUT_TEMPR93[17] ), .D(\A_DOUT_TEMPR94[17] ), .Y(
        OR4_128_Y));
    OR4 OR4_751 (.A(\A_DOUT_TEMPR8[34] ), .B(\A_DOUT_TEMPR9[34] ), .C(
        \A_DOUT_TEMPR10[34] ), .D(\A_DOUT_TEMPR11[34] ), .Y(OR4_751_Y));
    OR4 OR4_2813 (.A(OR4_2871_Y), .B(OR4_722_Y), .C(OR4_378_Y), .D(
        OR4_1877_Y), .Y(OR4_2813_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%37%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R37C7 (
        .A_DOUT({nc26370, nc26371, nc26372, nc26373, nc26374, nc26375, 
        nc26376, nc26377, nc26378, nc26379, nc26380, nc26381, nc26382, 
        nc26383, nc26384, \A_DOUT_TEMPR37[39] , \A_DOUT_TEMPR37[38] , 
        \A_DOUT_TEMPR37[37] , \A_DOUT_TEMPR37[36] , 
        \A_DOUT_TEMPR37[35] }), .B_DOUT({nc26385, nc26386, nc26387, 
        nc26388, nc26389, nc26390, nc26391, nc26392, nc26393, nc26394, 
        nc26395, nc26396, nc26397, nc26398, nc26399, 
        \B_DOUT_TEMPR37[39] , \B_DOUT_TEMPR37[38] , 
        \B_DOUT_TEMPR37[37] , \B_DOUT_TEMPR37[36] , 
        \B_DOUT_TEMPR37[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[37][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%64%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R64C2 (
        .A_DOUT({nc26400, nc26401, nc26402, nc26403, nc26404, nc26405, 
        nc26406, nc26407, nc26408, nc26409, nc26410, nc26411, nc26412, 
        nc26413, nc26414, \A_DOUT_TEMPR64[14] , \A_DOUT_TEMPR64[13] , 
        \A_DOUT_TEMPR64[12] , \A_DOUT_TEMPR64[11] , 
        \A_DOUT_TEMPR64[10] }), .B_DOUT({nc26415, nc26416, nc26417, 
        nc26418, nc26419, nc26420, nc26421, nc26422, nc26423, nc26424, 
        nc26425, nc26426, nc26427, nc26428, nc26429, 
        \B_DOUT_TEMPR64[14] , \B_DOUT_TEMPR64[13] , 
        \B_DOUT_TEMPR64[12] , \B_DOUT_TEMPR64[11] , 
        \B_DOUT_TEMPR64[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[64][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_348 (.A(OR4_2650_Y), .B(OR4_2964_Y), .C(OR4_2587_Y), .D(
        OR4_2977_Y), .Y(OR4_348_Y));
    OR4 OR4_329 (.A(\A_DOUT_TEMPR95[10] ), .B(\A_DOUT_TEMPR96[10] ), 
        .C(\A_DOUT_TEMPR97[10] ), .D(\A_DOUT_TEMPR98[10] ), .Y(
        OR4_329_Y));
    OR4 \OR4_B_DOUT[4]  (.A(OR4_925_Y), .B(OR4_121_Y), .C(OR4_1690_Y), 
        .D(OR4_2824_Y), .Y(B_DOUT[4]));
    OR4 OR4_2719 (.A(OR4_633_Y), .B(OR4_2122_Y), .C(OR4_2728_Y), .D(
        OR4_2518_Y), .Y(OR4_2719_Y));
    OR4 OR4_745 (.A(OR4_248_Y), .B(OR4_1196_Y), .C(OR4_827_Y), .D(
        OR4_2303_Y), .Y(OR4_745_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%28%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R28C2 (
        .A_DOUT({nc26430, nc26431, nc26432, nc26433, nc26434, nc26435, 
        nc26436, nc26437, nc26438, nc26439, nc26440, nc26441, nc26442, 
        nc26443, nc26444, \A_DOUT_TEMPR28[14] , \A_DOUT_TEMPR28[13] , 
        \A_DOUT_TEMPR28[12] , \A_DOUT_TEMPR28[11] , 
        \A_DOUT_TEMPR28[10] }), .B_DOUT({nc26445, nc26446, nc26447, 
        nc26448, nc26449, nc26450, nc26451, nc26452, nc26453, nc26454, 
        nc26455, nc26456, nc26457, nc26458, nc26459, 
        \B_DOUT_TEMPR28[14] , \B_DOUT_TEMPR28[13] , 
        \B_DOUT_TEMPR28[12] , \B_DOUT_TEMPR28[11] , 
        \B_DOUT_TEMPR28[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2268 (.A(\B_DOUT_TEMPR20[11] ), .B(\B_DOUT_TEMPR21[11] ), 
        .C(\B_DOUT_TEMPR22[11] ), .D(\B_DOUT_TEMPR23[11] ), .Y(
        OR4_2268_Y));
    OR4 OR4_986 (.A(\A_DOUT_TEMPR12[30] ), .B(\A_DOUT_TEMPR13[30] ), 
        .C(\A_DOUT_TEMPR14[30] ), .D(\A_DOUT_TEMPR15[30] ), .Y(
        OR4_986_Y));
    OR4 OR4_315 (.A(OR4_915_Y), .B(OR4_710_Y), .C(OR2_19_Y), .D(
        \A_DOUT_TEMPR74[39] ), .Y(OR4_315_Y));
    OR4 OR4_2592 (.A(\B_DOUT_TEMPR83[29] ), .B(\B_DOUT_TEMPR84[29] ), 
        .C(\B_DOUT_TEMPR85[29] ), .D(\B_DOUT_TEMPR86[29] ), .Y(
        OR4_2592_Y));
    OR4 OR4_2771 (.A(OR4_1637_Y), .B(OR4_2648_Y), .C(OR4_278_Y), .D(
        OR4_1952_Y), .Y(OR4_2771_Y));
    OR4 OR4_1410 (.A(\A_DOUT_TEMPR95[31] ), .B(\A_DOUT_TEMPR96[31] ), 
        .C(\A_DOUT_TEMPR97[31] ), .D(\A_DOUT_TEMPR98[31] ), .Y(
        OR4_1410_Y));
    OR2 OR2_65 (.A(\A_DOUT_TEMPR72[11] ), .B(\A_DOUT_TEMPR73[11] ), .Y(
        OR2_65_Y));
    OR4 OR4_839 (.A(OR4_1181_Y), .B(OR4_2846_Y), .C(OR4_2179_Y), .D(
        OR4_1527_Y), .Y(OR4_839_Y));
    OR4 OR4_707 (.A(OR4_2415_Y), .B(OR4_1442_Y), .C(OR4_1638_Y), .D(
        OR4_1452_Y), .Y(OR4_707_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%104%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R104C4 (
        .A_DOUT({nc26460, nc26461, nc26462, nc26463, nc26464, nc26465, 
        nc26466, nc26467, nc26468, nc26469, nc26470, nc26471, nc26472, 
        nc26473, nc26474, \A_DOUT_TEMPR104[24] , \A_DOUT_TEMPR104[23] , 
        \A_DOUT_TEMPR104[22] , \A_DOUT_TEMPR104[21] , 
        \A_DOUT_TEMPR104[20] }), .B_DOUT({nc26475, nc26476, nc26477, 
        nc26478, nc26479, nc26480, nc26481, nc26482, nc26483, nc26484, 
        nc26485, nc26486, nc26487, nc26488, nc26489, 
        \B_DOUT_TEMPR104[24] , \B_DOUT_TEMPR104[23] , 
        \B_DOUT_TEMPR104[22] , \B_DOUT_TEMPR104[21] , 
        \B_DOUT_TEMPR104[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[104][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_303 (.A(\B_DOUT_TEMPR52[19] ), .B(\B_DOUT_TEMPR53[19] ), 
        .C(\B_DOUT_TEMPR54[19] ), .D(\B_DOUT_TEMPR55[19] ), .Y(
        OR4_303_Y));
    OR4 OR4_852 (.A(\B_DOUT_TEMPR52[22] ), .B(\B_DOUT_TEMPR53[22] ), 
        .C(\B_DOUT_TEMPR54[22] ), .D(\B_DOUT_TEMPR55[22] ), .Y(
        OR4_852_Y));
    OR4 OR4_2116 (.A(\A_DOUT_TEMPR16[17] ), .B(\A_DOUT_TEMPR17[17] ), 
        .C(\A_DOUT_TEMPR18[17] ), .D(\A_DOUT_TEMPR19[17] ), .Y(
        OR4_2116_Y));
    OR4 OR4_2620 (.A(\B_DOUT_TEMPR103[29] ), .B(\B_DOUT_TEMPR104[29] ), 
        .C(\B_DOUT_TEMPR105[29] ), .D(\B_DOUT_TEMPR106[29] ), .Y(
        OR4_2620_Y));
    OR2 OR2_15 (.A(\A_DOUT_TEMPR72[28] ), .B(\A_DOUT_TEMPR73[28] ), .Y(
        OR2_15_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%47%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R47C1 (
        .A_DOUT({nc26490, nc26491, nc26492, nc26493, nc26494, nc26495, 
        nc26496, nc26497, nc26498, nc26499, nc26500, nc26501, nc26502, 
        nc26503, nc26504, \A_DOUT_TEMPR47[9] , \A_DOUT_TEMPR47[8] , 
        \A_DOUT_TEMPR47[7] , \A_DOUT_TEMPR47[6] , \A_DOUT_TEMPR47[5] })
        , .B_DOUT({nc26505, nc26506, nc26507, nc26508, nc26509, 
        nc26510, nc26511, nc26512, nc26513, nc26514, nc26515, nc26516, 
        nc26517, nc26518, nc26519, \B_DOUT_TEMPR47[9] , 
        \B_DOUT_TEMPR47[8] , \B_DOUT_TEMPR47[7] , \B_DOUT_TEMPR47[6] , 
        \B_DOUT_TEMPR47[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%63%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R63C7 (
        .A_DOUT({nc26520, nc26521, nc26522, nc26523, nc26524, nc26525, 
        nc26526, nc26527, nc26528, nc26529, nc26530, nc26531, nc26532, 
        nc26533, nc26534, \A_DOUT_TEMPR63[39] , \A_DOUT_TEMPR63[38] , 
        \A_DOUT_TEMPR63[37] , \A_DOUT_TEMPR63[36] , 
        \A_DOUT_TEMPR63[35] }), .B_DOUT({nc26535, nc26536, nc26537, 
        nc26538, nc26539, nc26540, nc26541, nc26542, nc26543, nc26544, 
        nc26545, nc26546, nc26547, nc26548, nc26549, 
        \B_DOUT_TEMPR63[39] , \B_DOUT_TEMPR63[38] , 
        \B_DOUT_TEMPR63[37] , \B_DOUT_TEMPR63[36] , 
        \B_DOUT_TEMPR63[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[63][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2518 (.A(\A_DOUT_TEMPR28[35] ), .B(\A_DOUT_TEMPR29[35] ), 
        .C(\A_DOUT_TEMPR30[35] ), .D(\A_DOUT_TEMPR31[35] ), .Y(
        OR4_2518_Y));
    OR4 OR4_708 (.A(\B_DOUT_TEMPR28[19] ), .B(\B_DOUT_TEMPR29[19] ), 
        .C(\B_DOUT_TEMPR30[19] ), .D(\B_DOUT_TEMPR31[19] ), .Y(
        OR4_708_Y));
    OR4 OR4_231 (.A(OR4_2903_Y), .B(OR4_1052_Y), .C(OR4_2076_Y), .D(
        OR4_76_Y), .Y(OR4_231_Y));
    OR2 OR2_4 (.A(\B_DOUT_TEMPR72[0] ), .B(\B_DOUT_TEMPR73[0] ), .Y(
        OR2_4_Y));
    OR4 OR4_831 (.A(OR4_1985_Y), .B(OR4_479_Y), .C(OR4_1131_Y), .D(
        OR4_291_Y), .Y(OR4_831_Y));
    OR4 OR4_1344 (.A(\A_DOUT_TEMPR36[9] ), .B(\A_DOUT_TEMPR37[9] ), .C(
        \A_DOUT_TEMPR38[9] ), .D(\A_DOUT_TEMPR39[9] ), .Y(OR4_1344_Y));
    OR4 OR4_2028 (.A(\B_DOUT_TEMPR12[34] ), .B(\B_DOUT_TEMPR13[34] ), 
        .C(\B_DOUT_TEMPR14[34] ), .D(\B_DOUT_TEMPR15[34] ), .Y(
        OR4_2028_Y));
    OR4 OR4_603 (.A(OR4_1560_Y), .B(OR4_2622_Y), .C(OR4_1293_Y), .D(
        OR4_2725_Y), .Y(OR4_603_Y));
    OR4 OR4_1184 (.A(\B_DOUT_TEMPR75[25] ), .B(\B_DOUT_TEMPR76[25] ), 
        .C(\B_DOUT_TEMPR77[25] ), .D(\B_DOUT_TEMPR78[25] ), .Y(
        OR4_1184_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%28%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R28C3 (
        .A_DOUT({nc26550, nc26551, nc26552, nc26553, nc26554, nc26555, 
        nc26556, nc26557, nc26558, nc26559, nc26560, nc26561, nc26562, 
        nc26563, nc26564, \A_DOUT_TEMPR28[19] , \A_DOUT_TEMPR28[18] , 
        \A_DOUT_TEMPR28[17] , \A_DOUT_TEMPR28[16] , 
        \A_DOUT_TEMPR28[15] }), .B_DOUT({nc26565, nc26566, nc26567, 
        nc26568, nc26569, nc26570, nc26571, nc26572, nc26573, nc26574, 
        nc26575, nc26576, nc26577, nc26578, nc26579, 
        \B_DOUT_TEMPR28[19] , \B_DOUT_TEMPR28[18] , 
        \B_DOUT_TEMPR28[17] , \B_DOUT_TEMPR28[16] , 
        \B_DOUT_TEMPR28[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[28][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_948 (.A(\A_DOUT_TEMPR40[27] ), .B(\A_DOUT_TEMPR41[27] ), 
        .C(\A_DOUT_TEMPR42[27] ), .D(\A_DOUT_TEMPR43[27] ), .Y(
        OR4_948_Y));
    OR4 OR4_1215 (.A(OR4_469_Y), .B(OR4_2034_Y), .C(OR4_2876_Y), .D(
        OR4_1888_Y), .Y(OR4_1215_Y));
    OR4 OR4_63 (.A(\B_DOUT_TEMPR44[20] ), .B(\B_DOUT_TEMPR45[20] ), .C(
        \B_DOUT_TEMPR46[20] ), .D(\B_DOUT_TEMPR47[20] ), .Y(OR4_63_Y));
    OR4 OR4_1751 (.A(\A_DOUT_TEMPR79[17] ), .B(\A_DOUT_TEMPR80[17] ), 
        .C(\A_DOUT_TEMPR81[17] ), .D(\A_DOUT_TEMPR82[17] ), .Y(
        OR4_1751_Y));
    OR4 OR4_222 (.A(OR4_2108_Y), .B(OR4_503_Y), .C(OR4_5_Y), .D(
        OR4_2601_Y), .Y(OR4_222_Y));
    OR4 OR4_2582 (.A(\A_DOUT_TEMPR44[9] ), .B(\A_DOUT_TEMPR45[9] ), .C(
        \A_DOUT_TEMPR46[9] ), .D(\A_DOUT_TEMPR47[9] ), .Y(OR4_2582_Y));
    OR4 OR4_199 (.A(\A_DOUT_TEMPR111[29] ), .B(\A_DOUT_TEMPR112[29] ), 
        .C(\A_DOUT_TEMPR113[29] ), .D(\A_DOUT_TEMPR114[29] ), .Y(
        OR4_199_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%24%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R24C1 (
        .A_DOUT({nc26580, nc26581, nc26582, nc26583, nc26584, nc26585, 
        nc26586, nc26587, nc26588, nc26589, nc26590, nc26591, nc26592, 
        nc26593, nc26594, \A_DOUT_TEMPR24[9] , \A_DOUT_TEMPR24[8] , 
        \A_DOUT_TEMPR24[7] , \A_DOUT_TEMPR24[6] , \A_DOUT_TEMPR24[5] })
        , .B_DOUT({nc26595, nc26596, nc26597, nc26598, nc26599, 
        nc26600, nc26601, nc26602, nc26603, nc26604, nc26605, nc26606, 
        nc26607, nc26608, nc26609, \B_DOUT_TEMPR24[9] , 
        \B_DOUT_TEMPR24[8] , \B_DOUT_TEMPR24[7] , \B_DOUT_TEMPR24[6] , 
        \B_DOUT_TEMPR24[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[24][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1290 (.A(\B_DOUT_TEMPR48[14] ), .B(\B_DOUT_TEMPR49[14] ), 
        .C(\B_DOUT_TEMPR50[14] ), .D(\B_DOUT_TEMPR51[14] ), .Y(
        OR4_1290_Y));
    OR4 \OR4_B_DOUT[11]  (.A(OR4_7_Y), .B(OR4_2599_Y), .C(OR4_908_Y), 
        .D(OR4_2928_Y), .Y(B_DOUT[11]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%20%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R20C4 (
        .A_DOUT({nc26610, nc26611, nc26612, nc26613, nc26614, nc26615, 
        nc26616, nc26617, nc26618, nc26619, nc26620, nc26621, nc26622, 
        nc26623, nc26624, \A_DOUT_TEMPR20[24] , \A_DOUT_TEMPR20[23] , 
        \A_DOUT_TEMPR20[22] , \A_DOUT_TEMPR20[21] , 
        \A_DOUT_TEMPR20[20] }), .B_DOUT({nc26625, nc26626, nc26627, 
        nc26628, nc26629, nc26630, nc26631, nc26632, nc26633, nc26634, 
        nc26635, nc26636, nc26637, nc26638, nc26639, 
        \B_DOUT_TEMPR20[24] , \B_DOUT_TEMPR20[23] , 
        \B_DOUT_TEMPR20[22] , \B_DOUT_TEMPR20[21] , 
        \B_DOUT_TEMPR20[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], B_DIN[22], 
        B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2450 (.A(\B_DOUT_TEMPR36[9] ), .B(\B_DOUT_TEMPR37[9] ), .C(
        \B_DOUT_TEMPR38[9] ), .D(\B_DOUT_TEMPR39[9] ), .Y(OR4_2450_Y));
    OR4 OR4_810 (.A(\A_DOUT_TEMPR68[12] ), .B(\A_DOUT_TEMPR69[12] ), 
        .C(\A_DOUT_TEMPR70[12] ), .D(\A_DOUT_TEMPR71[12] ), .Y(
        OR4_810_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%77%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R77C0 (
        .A_DOUT({nc26640, nc26641, nc26642, nc26643, nc26644, nc26645, 
        nc26646, nc26647, nc26648, nc26649, nc26650, nc26651, nc26652, 
        nc26653, nc26654, \A_DOUT_TEMPR77[4] , \A_DOUT_TEMPR77[3] , 
        \A_DOUT_TEMPR77[2] , \A_DOUT_TEMPR77[1] , \A_DOUT_TEMPR77[0] })
        , .B_DOUT({nc26655, nc26656, nc26657, nc26658, nc26659, 
        nc26660, nc26661, nc26662, nc26663, nc26664, nc26665, nc26666, 
        nc26667, nc26668, nc26669, \B_DOUT_TEMPR77[4] , 
        \B_DOUT_TEMPR77[3] , \B_DOUT_TEMPR77[2] , \B_DOUT_TEMPR77[1] , 
        \B_DOUT_TEMPR77[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[77][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1264 (.A(\A_DOUT_TEMPR48[14] ), .B(\A_DOUT_TEMPR49[14] ), 
        .C(\A_DOUT_TEMPR50[14] ), .D(\A_DOUT_TEMPR51[14] ), .Y(
        OR4_1264_Y));
    OR4 OR4_510 (.A(\B_DOUT_TEMPR0[23] ), .B(\B_DOUT_TEMPR1[23] ), .C(
        \B_DOUT_TEMPR2[23] ), .D(\B_DOUT_TEMPR3[23] ), .Y(OR4_510_Y));
    OR4 OR4_873 (.A(\B_DOUT_TEMPR0[11] ), .B(\B_DOUT_TEMPR1[11] ), .C(
        \B_DOUT_TEMPR2[11] ), .D(\B_DOUT_TEMPR3[11] ), .Y(OR4_873_Y));
    OR4 OR4_148 (.A(\A_DOUT_TEMPR111[30] ), .B(\A_DOUT_TEMPR112[30] ), 
        .C(\A_DOUT_TEMPR113[30] ), .D(\A_DOUT_TEMPR114[30] ), .Y(
        OR4_148_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%16%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R16C0 (
        .A_DOUT({nc26670, nc26671, nc26672, nc26673, nc26674, nc26675, 
        nc26676, nc26677, nc26678, nc26679, nc26680, nc26681, nc26682, 
        nc26683, nc26684, \A_DOUT_TEMPR16[4] , \A_DOUT_TEMPR16[3] , 
        \A_DOUT_TEMPR16[2] , \A_DOUT_TEMPR16[1] , \A_DOUT_TEMPR16[0] })
        , .B_DOUT({nc26685, nc26686, nc26687, nc26688, nc26689, 
        nc26690, nc26691, nc26692, nc26693, nc26694, nc26695, nc26696, 
        nc26697, nc26698, nc26699, \B_DOUT_TEMPR16[4] , 
        \B_DOUT_TEMPR16[3] , \B_DOUT_TEMPR16[2] , \B_DOUT_TEMPR16[1] , 
        \B_DOUT_TEMPR16[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[16][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2473 (.A(\A_DOUT_TEMPR52[11] ), .B(\A_DOUT_TEMPR53[11] ), 
        .C(\A_DOUT_TEMPR54[11] ), .D(\A_DOUT_TEMPR55[11] ), .Y(
        OR4_2473_Y));
    OR4 OR4_766 (.A(\B_DOUT_TEMPR52[28] ), .B(\B_DOUT_TEMPR53[28] ), 
        .C(\B_DOUT_TEMPR54[28] ), .D(\B_DOUT_TEMPR55[28] ), .Y(
        OR4_766_Y));
    OR4 OR4_349 (.A(OR4_638_Y), .B(OR4_1958_Y), .C(OR4_1595_Y), .D(
        OR4_2663_Y), .Y(OR4_349_Y));
    OR4 \OR4_A_DOUT[6]  (.A(OR4_1785_Y), .B(OR4_1343_Y), .C(OR4_2416_Y)
        , .D(OR4_2374_Y), .Y(A_DOUT[6]));
    OR4 OR4_1885 (.A(\A_DOUT_TEMPR115[39] ), .B(\A_DOUT_TEMPR116[39] ), 
        .C(\A_DOUT_TEMPR117[39] ), .D(\A_DOUT_TEMPR118[39] ), .Y(
        OR4_1885_Y));
    CFG1 #( .INIT(2'h1) )  \INVBLKX0[0]  (.A(A_ADDR[12]), .Y(
        \BLKX0[0] ));
    OR4 OR4_2255 (.A(\A_DOUT_TEMPR16[2] ), .B(\A_DOUT_TEMPR17[2] ), .C(
        \A_DOUT_TEMPR18[2] ), .D(\A_DOUT_TEMPR19[2] ), .Y(OR4_2255_Y));
    OR4 OR4_714 (.A(\A_DOUT_TEMPR40[3] ), .B(\A_DOUT_TEMPR41[3] ), .C(
        \A_DOUT_TEMPR42[3] ), .D(\A_DOUT_TEMPR43[3] ), .Y(OR4_714_Y));
    OR4 OR4_2090 (.A(\B_DOUT_TEMPR20[28] ), .B(\B_DOUT_TEMPR21[28] ), 
        .C(\B_DOUT_TEMPR22[28] ), .D(\B_DOUT_TEMPR23[28] ), .Y(
        OR4_2090_Y));
    OR4 OR4_1396 (.A(OR4_151_Y), .B(OR4_1711_Y), .C(OR4_2559_Y), .D(
        OR4_1581_Y), .Y(OR4_1396_Y));
    OR4 OR4_1063 (.A(\A_DOUT_TEMPR64[5] ), .B(\A_DOUT_TEMPR65[5] ), .C(
        \A_DOUT_TEMPR66[5] ), .D(\A_DOUT_TEMPR67[5] ), .Y(OR4_1063_Y));
    OR4 OR4_2124 (.A(OR4_1145_Y), .B(OR4_962_Y), .C(OR2_26_Y), .D(
        \B_DOUT_TEMPR74[30] ), .Y(OR4_2124_Y));
    OR4 \OR4_B_DOUT[12]  (.A(OR4_2959_Y), .B(OR4_696_Y), .C(OR4_2681_Y)
        , .D(OR4_2465_Y), .Y(B_DOUT[12]));
    OR4 OR4_1661 (.A(OR4_873_Y), .B(OR4_2408_Y), .C(OR4_198_Y), .D(
        OR4_2254_Y), .Y(OR4_1661_Y));
    OR4 OR4_337 (.A(\A_DOUT_TEMPR99[8] ), .B(\A_DOUT_TEMPR100[8] ), .C(
        \A_DOUT_TEMPR101[8] ), .D(\A_DOUT_TEMPR102[8] ), .Y(OR4_337_Y));
    OR4 OR4_1453 (.A(\B_DOUT_TEMPR8[13] ), .B(\B_DOUT_TEMPR9[13] ), .C(
        \B_DOUT_TEMPR10[13] ), .D(\B_DOUT_TEMPR11[13] ), .Y(OR4_1453_Y)
        );
    OR4 OR4_2808 (.A(OR4_2530_Y), .B(OR4_1847_Y), .C(OR4_724_Y), .D(
        OR4_1436_Y), .Y(OR4_2808_Y));
    OR4 OR4_1572 (.A(OR4_718_Y), .B(OR4_1538_Y), .C(OR4_602_Y), .D(
        OR4_2517_Y), .Y(OR4_1572_Y));
    OR4 OR4_3025 (.A(\A_DOUT_TEMPR16[11] ), .B(\A_DOUT_TEMPR17[11] ), 
        .C(\A_DOUT_TEMPR18[11] ), .D(\A_DOUT_TEMPR19[11] ), .Y(
        OR4_3025_Y));
    OR4 OR4_1763 (.A(\A_DOUT_TEMPR83[25] ), .B(\A_DOUT_TEMPR84[25] ), 
        .C(\A_DOUT_TEMPR85[25] ), .D(\A_DOUT_TEMPR86[25] ), .Y(
        OR4_1763_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%63%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R63C0 (
        .A_DOUT({nc26700, nc26701, nc26702, nc26703, nc26704, nc26705, 
        nc26706, nc26707, nc26708, nc26709, nc26710, nc26711, nc26712, 
        nc26713, nc26714, \A_DOUT_TEMPR63[4] , \A_DOUT_TEMPR63[3] , 
        \A_DOUT_TEMPR63[2] , \A_DOUT_TEMPR63[1] , \A_DOUT_TEMPR63[0] })
        , .B_DOUT({nc26715, nc26716, nc26717, nc26718, nc26719, 
        nc26720, nc26721, nc26722, nc26723, nc26724, nc26725, nc26726, 
        nc26727, nc26728, nc26729, \B_DOUT_TEMPR63[4] , 
        \B_DOUT_TEMPR63[3] , \B_DOUT_TEMPR63[2] , \B_DOUT_TEMPR63[1] , 
        \B_DOUT_TEMPR63[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[63][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_172 (.A(\A_DOUT_TEMPR40[15] ), .B(\A_DOUT_TEMPR41[15] ), 
        .C(\A_DOUT_TEMPR42[15] ), .D(\A_DOUT_TEMPR43[15] ), .Y(
        OR4_172_Y));
    OR4 OR4_838 (.A(OR4_2117_Y), .B(OR4_639_Y), .C(OR4_1350_Y), .D(
        OR4_1621_Y), .Y(OR4_838_Y));
    OR4 OR4_631 (.A(\B_DOUT_TEMPR83[24] ), .B(\B_DOUT_TEMPR84[24] ), 
        .C(\B_DOUT_TEMPR85[24] ), .D(\B_DOUT_TEMPR86[24] ), .Y(
        OR4_631_Y));
    OR4 OR4_1165 (.A(OR4_1044_Y), .B(OR4_1879_Y), .C(OR4_1080_Y), .D(
        OR4_6_Y), .Y(OR4_1165_Y));
    OR4 OR4_791 (.A(\B_DOUT_TEMPR75[31] ), .B(\B_DOUT_TEMPR76[31] ), 
        .C(\B_DOUT_TEMPR77[31] ), .D(\B_DOUT_TEMPR78[31] ), .Y(
        OR4_791_Y));
    OR4 OR4_917 (.A(\B_DOUT_TEMPR91[28] ), .B(\B_DOUT_TEMPR92[28] ), 
        .C(\B_DOUT_TEMPR93[28] ), .D(\B_DOUT_TEMPR94[28] ), .Y(
        OR4_917_Y));
    OR4 OR4_2645 (.A(\A_DOUT_TEMPR95[24] ), .B(\A_DOUT_TEMPR96[24] ), 
        .C(\A_DOUT_TEMPR97[24] ), .D(\A_DOUT_TEMPR98[24] ), .Y(
        OR4_2645_Y));
    OR4 OR4_561 (.A(\B_DOUT_TEMPR20[18] ), .B(\B_DOUT_TEMPR21[18] ), 
        .C(\B_DOUT_TEMPR22[18] ), .D(\B_DOUT_TEMPR23[18] ), .Y(
        OR4_561_Y));
    OR4 OR4_1907 (.A(\A_DOUT_TEMPR0[26] ), .B(\A_DOUT_TEMPR1[26] ), .C(
        \A_DOUT_TEMPR2[26] ), .D(\A_DOUT_TEMPR3[26] ), .Y(OR4_1907_Y));
    OR4 OR4_568 (.A(\B_DOUT_TEMPR64[34] ), .B(\B_DOUT_TEMPR65[34] ), 
        .C(\B_DOUT_TEMPR66[34] ), .D(\B_DOUT_TEMPR67[34] ), .Y(
        OR4_568_Y));
    OR4 OR4_2080 (.A(\B_DOUT_TEMPR32[15] ), .B(\B_DOUT_TEMPR33[15] ), 
        .C(\B_DOUT_TEMPR34[15] ), .D(\B_DOUT_TEMPR35[15] ), .Y(
        OR4_2080_Y));
    OR4 OR4_482 (.A(OR4_2314_Y), .B(OR4_102_Y), .C(OR2_50_Y), .D(
        \B_DOUT_TEMPR74[27] ), .Y(OR4_482_Y));
    OR4 OR4_242 (.A(\A_DOUT_TEMPR111[11] ), .B(\A_DOUT_TEMPR112[11] ), 
        .C(\A_DOUT_TEMPR113[11] ), .D(\A_DOUT_TEMPR114[11] ), .Y(
        OR4_242_Y));
    OR4 OR4_975 (.A(OR4_2190_Y), .B(OR4_1254_Y), .C(OR4_1441_Y), .D(
        OR4_1269_Y), .Y(OR4_975_Y));
    OR4 OR4_2514 (.A(\A_DOUT_TEMPR32[15] ), .B(\A_DOUT_TEMPR33[15] ), 
        .C(\A_DOUT_TEMPR34[15] ), .D(\A_DOUT_TEMPR35[15] ), .Y(
        OR4_2514_Y));
    OR4 OR4_2338 (.A(\B_DOUT_TEMPR68[28] ), .B(\B_DOUT_TEMPR69[28] ), 
        .C(\B_DOUT_TEMPR70[28] ), .D(\B_DOUT_TEMPR71[28] ), .Y(
        OR4_2338_Y));
    OR4 OR4_475 (.A(\B_DOUT_TEMPR83[19] ), .B(\B_DOUT_TEMPR84[19] ), 
        .C(\B_DOUT_TEMPR85[19] ), .D(\B_DOUT_TEMPR86[19] ), .Y(
        OR4_475_Y));
    OR4 OR4_803 (.A(\B_DOUT_TEMPR56[33] ), .B(\B_DOUT_TEMPR57[33] ), 
        .C(\B_DOUT_TEMPR58[33] ), .D(\B_DOUT_TEMPR59[33] ), .Y(
        OR4_803_Y));
    OR4 OR4_757 (.A(\B_DOUT_TEMPR79[37] ), .B(\B_DOUT_TEMPR80[37] ), 
        .C(\B_DOUT_TEMPR81[37] ), .D(\B_DOUT_TEMPR82[37] ), .Y(
        OR4_757_Y));
    OR4 OR4_43 (.A(\A_DOUT_TEMPR16[27] ), .B(\A_DOUT_TEMPR17[27] ), .C(
        \A_DOUT_TEMPR18[27] ), .D(\A_DOUT_TEMPR19[27] ), .Y(OR4_43_Y));
    OR4 OR4_1440 (.A(\B_DOUT_TEMPR79[24] ), .B(\B_DOUT_TEMPR80[24] ), 
        .C(\B_DOUT_TEMPR81[24] ), .D(\B_DOUT_TEMPR82[24] ), .Y(
        OR4_1440_Y));
    OR4 OR4_353 (.A(\B_DOUT_TEMPR32[4] ), .B(\B_DOUT_TEMPR33[4] ), .C(
        \B_DOUT_TEMPR34[4] ), .D(\B_DOUT_TEMPR35[4] ), .Y(OR4_353_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%67%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R67C7 (
        .A_DOUT({nc26730, nc26731, nc26732, nc26733, nc26734, nc26735, 
        nc26736, nc26737, nc26738, nc26739, nc26740, nc26741, nc26742, 
        nc26743, nc26744, \A_DOUT_TEMPR67[39] , \A_DOUT_TEMPR67[38] , 
        \A_DOUT_TEMPR67[37] , \A_DOUT_TEMPR67[36] , 
        \A_DOUT_TEMPR67[35] }), .B_DOUT({nc26745, nc26746, nc26747, 
        nc26748, nc26749, nc26750, nc26751, nc26752, nc26753, nc26754, 
        nc26755, nc26756, nc26757, nc26758, nc26759, 
        \B_DOUT_TEMPR67[39] , \B_DOUT_TEMPR67[38] , 
        \B_DOUT_TEMPR67[37] , \B_DOUT_TEMPR67[36] , 
        \B_DOUT_TEMPR67[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[67][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[16] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[16] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2825 (.A(\B_DOUT_TEMPR107[31] ), .B(\B_DOUT_TEMPR108[31] ), 
        .C(\B_DOUT_TEMPR109[31] ), .D(\B_DOUT_TEMPR110[31] ), .Y(
        OR4_2825_Y));
    OR4 OR4_1616 (.A(\A_DOUT_TEMPR83[14] ), .B(\A_DOUT_TEMPR84[14] ), 
        .C(\A_DOUT_TEMPR85[14] ), .D(\A_DOUT_TEMPR86[14] ), .Y(
        OR4_1616_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%14%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R14C2 (
        .A_DOUT({nc26760, nc26761, nc26762, nc26763, nc26764, nc26765, 
        nc26766, nc26767, nc26768, nc26769, nc26770, nc26771, nc26772, 
        nc26773, nc26774, \A_DOUT_TEMPR14[14] , \A_DOUT_TEMPR14[13] , 
        \A_DOUT_TEMPR14[12] , \A_DOUT_TEMPR14[11] , 
        \A_DOUT_TEMPR14[10] }), .B_DOUT({nc26775, nc26776, nc26777, 
        nc26778, nc26779, nc26780, nc26781, nc26782, nc26783, nc26784, 
        nc26785, nc26786, nc26787, nc26788, nc26789, 
        \B_DOUT_TEMPR14[14] , \B_DOUT_TEMPR14[13] , 
        \B_DOUT_TEMPR14[12] , \B_DOUT_TEMPR14[11] , 
        \B_DOUT_TEMPR14[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[14][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_434 (.A(\B_DOUT_TEMPR28[22] ), .B(\B_DOUT_TEMPR29[22] ), 
        .C(\B_DOUT_TEMPR30[22] ), .D(\B_DOUT_TEMPR31[22] ), .Y(
        OR4_434_Y));
    OR4 OR4_516 (.A(\B_DOUT_TEMPR32[33] ), .B(\B_DOUT_TEMPR33[33] ), 
        .C(\B_DOUT_TEMPR34[33] ), .D(\B_DOUT_TEMPR35[33] ), .Y(
        OR4_516_Y));
    OR4 OR4_1338 (.A(\A_DOUT_TEMPR56[5] ), .B(\A_DOUT_TEMPR57[5] ), .C(
        \A_DOUT_TEMPR58[5] ), .D(\A_DOUT_TEMPR59[5] ), .Y(OR4_1338_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%22%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R22C2 (
        .A_DOUT({nc26790, nc26791, nc26792, nc26793, nc26794, nc26795, 
        nc26796, nc26797, nc26798, nc26799, nc26800, nc26801, nc26802, 
        nc26803, nc26804, \A_DOUT_TEMPR22[14] , \A_DOUT_TEMPR22[13] , 
        \A_DOUT_TEMPR22[12] , \A_DOUT_TEMPR22[11] , 
        \A_DOUT_TEMPR22[10] }), .B_DOUT({nc26805, nc26806, nc26807, 
        nc26808, nc26809, nc26810, nc26811, nc26812, nc26813, nc26814, 
        nc26815, nc26816, nc26817, nc26818, nc26819, 
        \B_DOUT_TEMPR22[14] , \B_DOUT_TEMPR22[13] , 
        \B_DOUT_TEMPR22[12] , \B_DOUT_TEMPR22[11] , 
        \B_DOUT_TEMPR22[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR2 OR2_69 (.A(\B_DOUT_TEMPR72[13] ), .B(\B_DOUT_TEMPR73[13] ), .Y(
        OR2_69_Y));
    OR4 OR4_1061 (.A(\B_DOUT_TEMPR111[5] ), .B(\B_DOUT_TEMPR112[5] ), 
        .C(\B_DOUT_TEMPR113[5] ), .D(\B_DOUT_TEMPR114[5] ), .Y(
        OR4_1061_Y));
    OR4 OR4_758 (.A(\B_DOUT_TEMPR91[13] ), .B(\B_DOUT_TEMPR92[13] ), 
        .C(\B_DOUT_TEMPR93[13] ), .D(\B_DOUT_TEMPR94[13] ), .Y(
        OR4_758_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%6%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R6C2 (
        .A_DOUT({nc26820, nc26821, nc26822, nc26823, nc26824, nc26825, 
        nc26826, nc26827, nc26828, nc26829, nc26830, nc26831, nc26832, 
        nc26833, nc26834, \A_DOUT_TEMPR6[14] , \A_DOUT_TEMPR6[13] , 
        \A_DOUT_TEMPR6[12] , \A_DOUT_TEMPR6[11] , \A_DOUT_TEMPR6[10] })
        , .B_DOUT({nc26835, nc26836, nc26837, nc26838, nc26839, 
        nc26840, nc26841, nc26842, nc26843, nc26844, nc26845, nc26846, 
        nc26847, nc26848, nc26849, \B_DOUT_TEMPR6[14] , 
        \B_DOUT_TEMPR6[13] , \B_DOUT_TEMPR6[12] , \B_DOUT_TEMPR6[11] , 
        \B_DOUT_TEMPR6[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[6][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1110 (.A(\A_DOUT_TEMPR4[26] ), .B(\A_DOUT_TEMPR5[26] ), .C(
        \A_DOUT_TEMPR6[26] ), .D(\A_DOUT_TEMPR7[26] ), .Y(OR4_1110_Y));
    OR4 OR4_2496 (.A(\A_DOUT_TEMPR28[25] ), .B(\A_DOUT_TEMPR29[25] ), 
        .C(\A_DOUT_TEMPR30[25] ), .D(\A_DOUT_TEMPR31[25] ), .Y(
        OR4_2496_Y));
    OR4 OR4_653 (.A(OR4_1227_Y), .B(OR4_1493_Y), .C(OR4_64_Y), .D(
        OR4_1008_Y), .Y(OR4_653_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[29]  (.A(CFG3_1_Y), .B(
        CFG3_18_Y), .Y(\BLKX2[29] ));
    OR4 OR4_892 (.A(\A_DOUT_TEMPR115[31] ), .B(\A_DOUT_TEMPR116[31] ), 
        .C(\A_DOUT_TEMPR117[31] ), .D(\A_DOUT_TEMPR118[31] ), .Y(
        OR4_892_Y));
    OR2 OR2_19 (.A(\A_DOUT_TEMPR72[39] ), .B(\A_DOUT_TEMPR73[39] ), .Y(
        OR2_19_Y));
    OR4 OR4_2647 (.A(\B_DOUT_TEMPR99[12] ), .B(\B_DOUT_TEMPR100[12] ), 
        .C(\B_DOUT_TEMPR101[12] ), .D(\B_DOUT_TEMPR102[12] ), .Y(
        OR4_2647_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%83%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R83C3 (
        .A_DOUT({nc26850, nc26851, nc26852, nc26853, nc26854, nc26855, 
        nc26856, nc26857, nc26858, nc26859, nc26860, nc26861, nc26862, 
        nc26863, nc26864, \A_DOUT_TEMPR83[19] , \A_DOUT_TEMPR83[18] , 
        \A_DOUT_TEMPR83[17] , \A_DOUT_TEMPR83[16] , 
        \A_DOUT_TEMPR83[15] }), .B_DOUT({nc26865, nc26866, nc26867, 
        nc26868, nc26869, nc26870, nc26871, nc26872, nc26873, nc26874, 
        nc26875, nc26876, nc26877, nc26878, nc26879, 
        \B_DOUT_TEMPR83[19] , \B_DOUT_TEMPR83[18] , 
        \B_DOUT_TEMPR83[17] , \B_DOUT_TEMPR83[16] , 
        \B_DOUT_TEMPR83[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[83][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_365 (.A(\A_DOUT_TEMPR48[23] ), .B(\A_DOUT_TEMPR49[23] ), 
        .C(\A_DOUT_TEMPR50[23] ), .D(\A_DOUT_TEMPR51[23] ), .Y(
        OR4_365_Y));
    OR4 OR4_1245 (.A(\A_DOUT_TEMPR91[28] ), .B(\A_DOUT_TEMPR92[28] ), 
        .C(\A_DOUT_TEMPR93[28] ), .D(\A_DOUT_TEMPR94[28] ), .Y(
        OR4_1245_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%111%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R111C0 (
        .A_DOUT({nc26880, nc26881, nc26882, nc26883, nc26884, nc26885, 
        nc26886, nc26887, nc26888, nc26889, nc26890, nc26891, nc26892, 
        nc26893, nc26894, \A_DOUT_TEMPR111[4] , \A_DOUT_TEMPR111[3] , 
        \A_DOUT_TEMPR111[2] , \A_DOUT_TEMPR111[1] , 
        \A_DOUT_TEMPR111[0] }), .B_DOUT({nc26895, nc26896, nc26897, 
        nc26898, nc26899, nc26900, nc26901, nc26902, nc26903, nc26904, 
        nc26905, nc26906, nc26907, nc26908, nc26909, 
        \B_DOUT_TEMPR111[4] , \B_DOUT_TEMPR111[3] , 
        \B_DOUT_TEMPR111[2] , \B_DOUT_TEMPR111[1] , 
        \B_DOUT_TEMPR111[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[111][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%85%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R85C3 (
        .A_DOUT({nc26910, nc26911, nc26912, nc26913, nc26914, nc26915, 
        nc26916, nc26917, nc26918, nc26919, nc26920, nc26921, nc26922, 
        nc26923, nc26924, \A_DOUT_TEMPR85[19] , \A_DOUT_TEMPR85[18] , 
        \A_DOUT_TEMPR85[17] , \A_DOUT_TEMPR85[16] , 
        \A_DOUT_TEMPR85[15] }), .B_DOUT({nc26925, nc26926, nc26927, 
        nc26928, nc26929, nc26930, nc26931, nc26932, nc26933, nc26934, 
        nc26935, nc26936, nc26937, nc26938, nc26939, 
        \B_DOUT_TEMPR85[19] , \B_DOUT_TEMPR85[18] , 
        \B_DOUT_TEMPR85[17] , \B_DOUT_TEMPR85[16] , 
        \B_DOUT_TEMPR85[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[85][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1800 (.A(\A_DOUT_TEMPR83[38] ), .B(\A_DOUT_TEMPR84[38] ), 
        .C(\A_DOUT_TEMPR85[38] ), .D(\A_DOUT_TEMPR86[38] ), .Y(
        OR4_1800_Y));
    OR4 OR4_1492 (.A(\B_DOUT_TEMPR111[14] ), .B(\B_DOUT_TEMPR112[14] ), 
        .C(\B_DOUT_TEMPR113[14] ), .D(\B_DOUT_TEMPR114[14] ), .Y(
        OR4_1492_Y));
    OR4 OR4_102 (.A(\B_DOUT_TEMPR68[27] ), .B(\B_DOUT_TEMPR69[27] ), 
        .C(\B_DOUT_TEMPR70[27] ), .D(\B_DOUT_TEMPR71[27] ), .Y(
        OR4_102_Y));
    OR4 \OR4_A_DOUT[30]  (.A(OR4_1571_Y), .B(OR4_824_Y), .C(OR4_1024_Y)
        , .D(OR4_2355_Y), .Y(A_DOUT[30]));
    OR4 OR4_2708 (.A(\B_DOUT_TEMPR91[16] ), .B(\B_DOUT_TEMPR92[16] ), 
        .C(\B_DOUT_TEMPR93[16] ), .D(\B_DOUT_TEMPR94[16] ), .Y(
        OR4_2708_Y));
    OR4 OR4_1498 (.A(\A_DOUT_TEMPR79[24] ), .B(\A_DOUT_TEMPR80[24] ), 
        .C(\A_DOUT_TEMPR81[24] ), .D(\A_DOUT_TEMPR82[24] ), .Y(
        OR4_1498_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%13%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R13C7 (
        .A_DOUT({nc26940, nc26941, nc26942, nc26943, nc26944, nc26945, 
        nc26946, nc26947, nc26948, nc26949, nc26950, nc26951, nc26952, 
        nc26953, nc26954, \A_DOUT_TEMPR13[39] , \A_DOUT_TEMPR13[38] , 
        \A_DOUT_TEMPR13[37] , \A_DOUT_TEMPR13[36] , 
        \A_DOUT_TEMPR13[35] }), .B_DOUT({nc26955, nc26956, nc26957, 
        nc26958, nc26959, nc26960, nc26961, nc26962, nc26963, nc26964, 
        nc26965, nc26966, nc26967, nc26968, nc26969, 
        \B_DOUT_TEMPR13[39] , \B_DOUT_TEMPR13[38] , 
        \B_DOUT_TEMPR13[37] , \B_DOUT_TEMPR13[36] , 
        \B_DOUT_TEMPR13[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2211 (.A(\A_DOUT_TEMPR111[2] ), .B(\A_DOUT_TEMPR112[2] ), 
        .C(\A_DOUT_TEMPR113[2] ), .D(\A_DOUT_TEMPR114[2] ), .Y(
        OR4_2211_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%91%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R91C5 (
        .A_DOUT({nc26970, nc26971, nc26972, nc26973, nc26974, nc26975, 
        nc26976, nc26977, nc26978, nc26979, nc26980, nc26981, nc26982, 
        nc26983, nc26984, \A_DOUT_TEMPR91[29] , \A_DOUT_TEMPR91[28] , 
        \A_DOUT_TEMPR91[27] , \A_DOUT_TEMPR91[26] , 
        \A_DOUT_TEMPR91[25] }), .B_DOUT({nc26985, nc26986, nc26987, 
        nc26988, nc26989, nc26990, nc26991, nc26992, nc26993, nc26994, 
        nc26995, nc26996, nc26997, nc26998, nc26999, 
        \B_DOUT_TEMPR91[29] , \B_DOUT_TEMPR91[28] , 
        \B_DOUT_TEMPR91[27] , \B_DOUT_TEMPR91[26] , 
        \B_DOUT_TEMPR91[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[91][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2795 (.A(\B_DOUT_TEMPR75[12] ), .B(\B_DOUT_TEMPR76[12] ), 
        .C(\B_DOUT_TEMPR77[12] ), .D(\B_DOUT_TEMPR78[12] ), .Y(
        OR4_2795_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%23%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R23C1 (
        .A_DOUT({nc27000, nc27001, nc27002, nc27003, nc27004, nc27005, 
        nc27006, nc27007, nc27008, nc27009, nc27010, nc27011, nc27012, 
        nc27013, nc27014, \A_DOUT_TEMPR23[9] , \A_DOUT_TEMPR23[8] , 
        \A_DOUT_TEMPR23[7] , \A_DOUT_TEMPR23[6] , \A_DOUT_TEMPR23[5] })
        , .B_DOUT({nc27015, nc27016, nc27017, nc27018, nc27019, 
        nc27020, nc27021, nc27022, nc27023, nc27024, nc27025, nc27026, 
        nc27027, nc27028, nc27029, \B_DOUT_TEMPR23[9] , 
        \B_DOUT_TEMPR23[8] , \B_DOUT_TEMPR23[7] , \B_DOUT_TEMPR23[6] , 
        \B_DOUT_TEMPR23[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[23][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], B_DIN[7], 
        B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[2] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_1070 (.A(OR4_665_Y), .B(OR4_984_Y), .C(OR4_596_Y), .D(
        OR4_1006_Y), .Y(OR4_1070_Y));
    OR4 OR4_2656 (.A(\B_DOUT_TEMPR32[23] ), .B(\B_DOUT_TEMPR33[23] ), 
        .C(\B_DOUT_TEMPR34[23] ), .D(\B_DOUT_TEMPR35[23] ), .Y(
        OR4_2656_Y));
    OR4 OR4_1804 (.A(\A_DOUT_TEMPR103[25] ), .B(\A_DOUT_TEMPR104[25] ), 
        .C(\A_DOUT_TEMPR105[25] ), .D(\A_DOUT_TEMPR106[25] ), .Y(
        OR4_1804_Y));
    OR4 OR4_2486 (.A(\A_DOUT_TEMPR60[11] ), .B(\A_DOUT_TEMPR61[11] ), 
        .C(\A_DOUT_TEMPR62[11] ), .D(\A_DOUT_TEMPR63[11] ), .Y(
        OR4_2486_Y));
    OR4 OR4_2150 (.A(\B_DOUT_TEMPR52[31] ), .B(\B_DOUT_TEMPR53[31] ), 
        .C(\B_DOUT_TEMPR54[31] ), .D(\B_DOUT_TEMPR55[31] ), .Y(
        OR4_2150_Y));
    OR4 OR4_905 (.A(\B_DOUT_TEMPR24[0] ), .B(\B_DOUT_TEMPR25[0] ), .C(
        \B_DOUT_TEMPR26[0] ), .D(\B_DOUT_TEMPR27[0] ), .Y(OR4_905_Y));
    OR4 OR4_405 (.A(\A_DOUT_TEMPR12[9] ), .B(\A_DOUT_TEMPR13[9] ), .C(
        \A_DOUT_TEMPR14[9] ), .D(\A_DOUT_TEMPR15[9] ), .Y(OR4_405_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%79%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R79C6 (
        .A_DOUT({nc27030, nc27031, nc27032, nc27033, nc27034, nc27035, 
        nc27036, nc27037, nc27038, nc27039, nc27040, nc27041, nc27042, 
        nc27043, nc27044, \A_DOUT_TEMPR79[34] , \A_DOUT_TEMPR79[33] , 
        \A_DOUT_TEMPR79[32] , \A_DOUT_TEMPR79[31] , 
        \A_DOUT_TEMPR79[30] }), .B_DOUT({nc27045, nc27046, nc27047, 
        nc27048, nc27049, nc27050, nc27051, nc27052, nc27053, nc27054, 
        nc27055, nc27056, nc27057, nc27058, nc27059, 
        \B_DOUT_TEMPR79[34] , \B_DOUT_TEMPR79[33] , 
        \B_DOUT_TEMPR79[32] , \B_DOUT_TEMPR79[31] , 
        \B_DOUT_TEMPR79[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[79][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2276 (.A(OR4_2148_Y), .B(OR4_735_Y), .C(OR4_300_Y), .D(
        OR4_1991_Y), .Y(OR4_2276_Y));
    OR4 OR4_2435 (.A(\B_DOUT_TEMPR111[38] ), .B(\B_DOUT_TEMPR112[38] ), 
        .C(\B_DOUT_TEMPR113[38] ), .D(\B_DOUT_TEMPR114[38] ), .Y(
        OR4_2435_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%41%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R41C0 (
        .A_DOUT({nc27060, nc27061, nc27062, nc27063, nc27064, nc27065, 
        nc27066, nc27067, nc27068, nc27069, nc27070, nc27071, nc27072, 
        nc27073, nc27074, \A_DOUT_TEMPR41[4] , \A_DOUT_TEMPR41[3] , 
        \A_DOUT_TEMPR41[2] , \A_DOUT_TEMPR41[1] , \A_DOUT_TEMPR41[0] })
        , .B_DOUT({nc27075, nc27076, nc27077, nc27078, nc27079, 
        nc27080, nc27081, nc27082, nc27083, nc27084, nc27085, nc27086, 
        nc27087, nc27088, nc27089, \B_DOUT_TEMPR41[4] , 
        \B_DOUT_TEMPR41[3] , \B_DOUT_TEMPR41[2] , \B_DOUT_TEMPR41[1] , 
        \B_DOUT_TEMPR41[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[41][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2562 (.A(\A_DOUT_TEMPR68[31] ), .B(\A_DOUT_TEMPR69[31] ), 
        .C(\A_DOUT_TEMPR70[31] ), .D(\A_DOUT_TEMPR71[31] ), .Y(
        OR4_2562_Y));
    OR4 OR4_1590 (.A(\B_DOUT_TEMPR20[16] ), .B(\B_DOUT_TEMPR21[16] ), 
        .C(\B_DOUT_TEMPR22[16] ), .D(\B_DOUT_TEMPR23[16] ), .Y(
        OR4_1590_Y));
    OR4 OR4_860 (.A(\B_DOUT_TEMPR40[16] ), .B(\B_DOUT_TEMPR41[16] ), 
        .C(\B_DOUT_TEMPR42[16] ), .D(\B_DOUT_TEMPR43[16] ), .Y(
        OR4_860_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%80%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R80C1 (
        .A_DOUT({nc27090, nc27091, nc27092, nc27093, nc27094, nc27095, 
        nc27096, nc27097, nc27098, nc27099, nc27100, nc27101, nc27102, 
        nc27103, nc27104, \A_DOUT_TEMPR80[9] , \A_DOUT_TEMPR80[8] , 
        \A_DOUT_TEMPR80[7] , \A_DOUT_TEMPR80[6] , \A_DOUT_TEMPR80[5] })
        , .B_DOUT({nc27105, nc27106, nc27107, nc27108, nc27109, 
        nc27110, nc27111, nc27112, nc27113, nc27114, nc27115, nc27116, 
        nc27117, nc27118, nc27119, \B_DOUT_TEMPR80[9] , 
        \B_DOUT_TEMPR80[8] , \B_DOUT_TEMPR80[7] , \B_DOUT_TEMPR80[6] , 
        \B_DOUT_TEMPR80[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[80][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1435 (.A(\A_DOUT_TEMPR8[39] ), .B(\A_DOUT_TEMPR9[39] ), .C(
        \A_DOUT_TEMPR10[39] ), .D(\A_DOUT_TEMPR11[39] ), .Y(OR4_1435_Y)
        );
    OR4 \OR4_B_DOUT[19]  (.A(OR4_641_Y), .B(OR4_1983_Y), .C(OR4_634_Y), 
        .D(OR4_2487_Y), .Y(B_DOUT[19]));
    OR4 OR4_560 (.A(OR4_2926_Y), .B(OR4_2731_Y), .C(OR4_2667_Y), .D(
        OR4_1483_Y), .Y(OR4_560_Y));
    OR4 OR4_2785 (.A(\B_DOUT_TEMPR75[29] ), .B(\B_DOUT_TEMPR76[29] ), 
        .C(\B_DOUT_TEMPR77[29] ), .D(\B_DOUT_TEMPR78[29] ), .Y(
        OR4_2785_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%3%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R3C6 (
        .A_DOUT({nc27120, nc27121, nc27122, nc27123, nc27124, nc27125, 
        nc27126, nc27127, nc27128, nc27129, nc27130, nc27131, nc27132, 
        nc27133, nc27134, \A_DOUT_TEMPR3[34] , \A_DOUT_TEMPR3[33] , 
        \A_DOUT_TEMPR3[32] , \A_DOUT_TEMPR3[31] , \A_DOUT_TEMPR3[30] })
        , .B_DOUT({nc27135, nc27136, nc27137, nc27138, nc27139, 
        nc27140, nc27141, nc27142, nc27143, nc27144, nc27145, nc27146, 
        nc27147, nc27148, nc27149, \B_DOUT_TEMPR3[34] , 
        \B_DOUT_TEMPR3[33] , \B_DOUT_TEMPR3[32] , \B_DOUT_TEMPR3[31] , 
        \B_DOUT_TEMPR3[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[3][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1256 (.A(OR4_1039_Y), .B(OR4_2183_Y), .C(OR4_201_Y), .D(
        OR4_2569_Y), .Y(OR4_1256_Y));
    OR4 OR4_1688 (.A(\A_DOUT_TEMPR107[0] ), .B(\A_DOUT_TEMPR108[0] ), 
        .C(\A_DOUT_TEMPR109[0] ), .D(\A_DOUT_TEMPR110[0] ), .Y(
        OR4_1688_Y));
    OR4 OR4_764 (.A(\A_DOUT_TEMPR12[19] ), .B(\A_DOUT_TEMPR13[19] ), 
        .C(\A_DOUT_TEMPR14[19] ), .D(\A_DOUT_TEMPR15[19] ), .Y(
        OR4_764_Y));
    OR4 OR4_2344 (.A(\B_DOUT_TEMPR32[11] ), .B(\B_DOUT_TEMPR33[11] ), 
        .C(\B_DOUT_TEMPR34[11] ), .D(\B_DOUT_TEMPR35[11] ), .Y(
        OR4_2344_Y));
    OR4 OR4_2736 (.A(\A_DOUT_TEMPR40[4] ), .B(\A_DOUT_TEMPR41[4] ), .C(
        \A_DOUT_TEMPR42[4] ), .D(\A_DOUT_TEMPR43[4] ), .Y(OR4_2736_Y));
    OR4 OR4_1476 (.A(OR4_2680_Y), .B(OR4_545_Y), .C(OR4_177_Y), .D(
        OR4_1677_Y), .Y(OR4_1476_Y));
    OR4 OR4_853 (.A(\A_DOUT_TEMPR44[32] ), .B(\A_DOUT_TEMPR45[32] ), 
        .C(\A_DOUT_TEMPR46[32] ), .D(\A_DOUT_TEMPR47[32] ), .Y(
        OR4_853_Y));
    OR4 OR4_834 (.A(\B_DOUT_TEMPR20[30] ), .B(\B_DOUT_TEMPR21[30] ), 
        .C(\B_DOUT_TEMPR22[30] ), .D(\B_DOUT_TEMPR23[30] ), .Y(
        OR4_834_Y));
    OR4 OR4_1913 (.A(OR4_507_Y), .B(OR4_2573_Y), .C(OR4_2797_Y), .D(
        OR4_2589_Y), .Y(OR4_1913_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%110%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R110C2 (
        .A_DOUT({nc27150, nc27151, nc27152, nc27153, nc27154, nc27155, 
        nc27156, nc27157, nc27158, nc27159, nc27160, nc27161, nc27162, 
        nc27163, nc27164, \A_DOUT_TEMPR110[14] , \A_DOUT_TEMPR110[13] , 
        \A_DOUT_TEMPR110[12] , \A_DOUT_TEMPR110[11] , 
        \A_DOUT_TEMPR110[10] }), .B_DOUT({nc27165, nc27166, nc27167, 
        nc27168, nc27169, nc27170, nc27171, nc27172, nc27173, nc27174, 
        nc27175, nc27176, nc27177, nc27178, nc27179, 
        \B_DOUT_TEMPR110[14] , \B_DOUT_TEMPR110[13] , 
        \B_DOUT_TEMPR110[12] , \B_DOUT_TEMPR110[11] , 
        \B_DOUT_TEMPR110[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[110][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1736 (.A(\A_DOUT_TEMPR44[15] ), .B(\A_DOUT_TEMPR45[15] ), 
        .C(\A_DOUT_TEMPR46[15] ), .D(\A_DOUT_TEMPR47[15] ), .Y(
        OR4_1736_Y));
    OR4 OR4_532 (.A(\B_DOUT_TEMPR103[2] ), .B(\B_DOUT_TEMPR104[2] ), 
        .C(\B_DOUT_TEMPR105[2] ), .D(\B_DOUT_TEMPR106[2] ), .Y(
        OR4_532_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%77%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R77C1 (
        .A_DOUT({nc27180, nc27181, nc27182, nc27183, nc27184, nc27185, 
        nc27186, nc27187, nc27188, nc27189, nc27190, nc27191, nc27192, 
        nc27193, nc27194, \A_DOUT_TEMPR77[9] , \A_DOUT_TEMPR77[8] , 
        \A_DOUT_TEMPR77[7] , \A_DOUT_TEMPR77[6] , \A_DOUT_TEMPR77[5] })
        , .B_DOUT({nc27195, nc27196, nc27197, nc27198, nc27199, 
        nc27200, nc27201, nc27202, nc27203, nc27204, nc27205, nc27206, 
        nc27207, nc27208, nc27209, \B_DOUT_TEMPR77[9] , 
        \B_DOUT_TEMPR77[8] , \B_DOUT_TEMPR77[7] , \B_DOUT_TEMPR77[6] , 
        \B_DOUT_TEMPR77[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[77][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%13%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R13C0 (
        .A_DOUT({nc27210, nc27211, nc27212, nc27213, nc27214, nc27215, 
        nc27216, nc27217, nc27218, nc27219, nc27220, nc27221, nc27222, 
        nc27223, nc27224, \A_DOUT_TEMPR13[4] , \A_DOUT_TEMPR13[3] , 
        \A_DOUT_TEMPR13[2] , \A_DOUT_TEMPR13[1] , \A_DOUT_TEMPR13[0] })
        , .B_DOUT({nc27225, nc27226, nc27227, nc27228, nc27229, 
        nc27230, nc27231, nc27232, nc27233, nc27234, nc27235, nc27236, 
        nc27237, nc27238, nc27239, \B_DOUT_TEMPR13[4] , 
        \B_DOUT_TEMPR13[3] , \B_DOUT_TEMPR13[2] , \B_DOUT_TEMPR13[1] , 
        \B_DOUT_TEMPR13[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[13][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[3] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    OR4 OR4_2876 (.A(\A_DOUT_TEMPR8[16] ), .B(\A_DOUT_TEMPR9[16] ), .C(
        \A_DOUT_TEMPR10[16] ), .D(\A_DOUT_TEMPR11[16] ), .Y(OR4_2876_Y)
        );
    OR4 OR4_1646 (.A(\B_DOUT_TEMPR8[24] ), .B(\B_DOUT_TEMPR9[24] ), .C(
        \B_DOUT_TEMPR10[24] ), .D(\B_DOUT_TEMPR11[24] ), .Y(OR4_1646_Y)
        );
    OR4 OR4_797 (.A(\A_DOUT_TEMPR32[39] ), .B(\A_DOUT_TEMPR33[39] ), 
        .C(\A_DOUT_TEMPR34[39] ), .D(\A_DOUT_TEMPR35[39] ), .Y(
        OR4_797_Y));
    OR4 OR4_1140 (.A(\B_DOUT_TEMPR40[32] ), .B(\B_DOUT_TEMPR41[32] ), 
        .C(\B_DOUT_TEMPR42[32] ), .D(\B_DOUT_TEMPR43[32] ), .Y(
        OR4_1140_Y));
    OR4 OR4_393 (.A(\B_DOUT_TEMPR44[3] ), .B(\B_DOUT_TEMPR45[3] ), .C(
        \B_DOUT_TEMPR46[3] ), .D(\B_DOUT_TEMPR47[3] ), .Y(OR4_393_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%8%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R8C2 (
        .A_DOUT({nc27240, nc27241, nc27242, nc27243, nc27244, nc27245, 
        nc27246, nc27247, nc27248, nc27249, nc27250, nc27251, nc27252, 
        nc27253, nc27254, \A_DOUT_TEMPR8[14] , \A_DOUT_TEMPR8[13] , 
        \A_DOUT_TEMPR8[12] , \A_DOUT_TEMPR8[11] , \A_DOUT_TEMPR8[10] })
        , .B_DOUT({nc27255, nc27256, nc27257, nc27258, nc27259, 
        nc27260, nc27261, nc27262, nc27263, nc27264, nc27265, nc27266, 
        nc27267, nc27268, nc27269, \B_DOUT_TEMPR8[14] , 
        \B_DOUT_TEMPR8[13] , \B_DOUT_TEMPR8[12] , \B_DOUT_TEMPR8[11] , 
        \B_DOUT_TEMPR8[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[8][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1995 (.A(\A_DOUT_TEMPR32[17] ), .B(\A_DOUT_TEMPR33[17] ), 
        .C(\A_DOUT_TEMPR34[17] ), .D(\A_DOUT_TEMPR35[17] ), .Y(
        OR4_1995_Y));
    OR4 OR4_967 (.A(OR4_2068_Y), .B(OR4_1104_Y), .C(OR4_1306_Y), .D(
        OR4_1117_Y), .Y(OR4_967_Y));
    OR4 OR4_1775 (.A(\B_DOUT_TEMPR83[31] ), .B(\B_DOUT_TEMPR84[31] ), 
        .C(\B_DOUT_TEMPR85[31] ), .D(\B_DOUT_TEMPR86[31] ), .Y(
        OR4_1775_Y));
    OR4 OR4_798 (.A(\B_DOUT_TEMPR91[0] ), .B(\B_DOUT_TEMPR92[0] ), .C(
        \B_DOUT_TEMPR93[0] ), .D(\B_DOUT_TEMPR94[0] ), .Y(OR4_798_Y));
    OR4 OR4_1311 (.A(\A_DOUT_TEMPR48[39] ), .B(\A_DOUT_TEMPR49[39] ), 
        .C(\A_DOUT_TEMPR50[39] ), .D(\A_DOUT_TEMPR51[39] ), .Y(
        OR4_1311_Y));
    OR4 OR4_97 (.A(\A_DOUT_TEMPR115[38] ), .B(\A_DOUT_TEMPR116[38] ), 
        .C(\A_DOUT_TEMPR117[38] ), .D(\A_DOUT_TEMPR118[38] ), .Y(
        OR4_97_Y));
    OR4 OR4_693 (.A(\B_DOUT_TEMPR4[9] ), .B(\B_DOUT_TEMPR5[9] ), .C(
        \B_DOUT_TEMPR6[9] ), .D(\B_DOUT_TEMPR7[9] ), .Y(OR4_693_Y));
    OR4 OR4_2060 (.A(OR4_760_Y), .B(OR4_1090_Y), .C(OR4_2686_Y), .D(
        OR4_550_Y), .Y(OR4_2060_Y));
    OR4 OR4_1699 (.A(\A_DOUT_TEMPR0[14] ), .B(\A_DOUT_TEMPR1[14] ), .C(
        \A_DOUT_TEMPR2[14] ), .D(\A_DOUT_TEMPR3[14] ), .Y(OR4_1699_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%17%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R17C7 (
        .A_DOUT({nc27270, nc27271, nc27272, nc27273, nc27274, nc27275, 
        nc27276, nc27277, nc27278, nc27279, nc27280, nc27281, nc27282, 
        nc27283, nc27284, \A_DOUT_TEMPR17[39] , \A_DOUT_TEMPR17[38] , 
        \A_DOUT_TEMPR17[37] , \A_DOUT_TEMPR17[36] , 
        \A_DOUT_TEMPR17[35] }), .B_DOUT({nc27285, nc27286, nc27287, 
        nc27288, nc27289, nc27290, nc27291, nc27292, nc27293, nc27294, 
        nc27295, nc27296, nc27297, nc27298, nc27299, 
        \B_DOUT_TEMPR17[39] , \B_DOUT_TEMPR17[38] , 
        \B_DOUT_TEMPR17[37] , \B_DOUT_TEMPR17[36] , 
        \B_DOUT_TEMPR17[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[17][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[4] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], B_DIN[37], 
        B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1856 (.A(OR4_2956_Y), .B(OR4_812_Y), .C(OR4_458_Y), .D(
        OR4_1957_Y), .Y(OR4_1856_Y));
    OR4 OR4_1811 (.A(\B_DOUT_TEMPR115[19] ), .B(\B_DOUT_TEMPR116[19] ), 
        .C(\B_DOUT_TEMPR117[19] ), .D(\B_DOUT_TEMPR118[19] ), .Y(
        OR4_1811_Y));
    OR4 OR4_152 (.A(\A_DOUT_TEMPR32[14] ), .B(\A_DOUT_TEMPR33[14] ), 
        .C(\A_DOUT_TEMPR34[14] ), .D(\A_DOUT_TEMPR35[14] ), .Y(
        OR4_152_Y));
    OR4 OR4_2953 (.A(\B_DOUT_TEMPR87[20] ), .B(\B_DOUT_TEMPR88[20] ), 
        .C(\B_DOUT_TEMPR89[20] ), .D(\B_DOUT_TEMPR90[20] ), .Y(
        OR4_2953_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%1%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R1C2 (
        .A_DOUT({nc27300, nc27301, nc27302, nc27303, nc27304, nc27305, 
        nc27306, nc27307, nc27308, nc27309, nc27310, nc27311, nc27312, 
        nc27313, nc27314, \A_DOUT_TEMPR1[14] , \A_DOUT_TEMPR1[13] , 
        \A_DOUT_TEMPR1[12] , \A_DOUT_TEMPR1[11] , \A_DOUT_TEMPR1[10] })
        , .B_DOUT({nc27315, nc27316, nc27317, nc27318, nc27319, 
        nc27320, nc27321, nc27322, nc27323, nc27324, nc27325, nc27326, 
        nc27327, nc27328, nc27329, \B_DOUT_TEMPR1[14] , 
        \B_DOUT_TEMPR1[13] , \B_DOUT_TEMPR1[12] , \B_DOUT_TEMPR1[11] , 
        \B_DOUT_TEMPR1[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[1][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[0] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_926 (.A(\A_DOUT_TEMPR32[12] ), .B(\A_DOUT_TEMPR33[12] ), 
        .C(\A_DOUT_TEMPR34[12] ), .D(\A_DOUT_TEMPR35[12] ), .Y(
        OR4_926_Y));
    OR4 OR4_566 (.A(\B_DOUT_TEMPR28[33] ), .B(\B_DOUT_TEMPR29[33] ), 
        .C(\B_DOUT_TEMPR30[33] ), .D(\B_DOUT_TEMPR31[33] ), .Y(
        OR4_566_Y));
    OR4 OR4_2628 (.A(OR4_2296_Y), .B(OR4_1333_Y), .C(OR4_2249_Y), .D(
        OR4_437_Y), .Y(OR4_2628_Y));
    OR4 OR4_2596 (.A(\A_DOUT_TEMPR48[15] ), .B(\A_DOUT_TEMPR49[15] ), 
        .C(\A_DOUT_TEMPR50[15] ), .D(\A_DOUT_TEMPR51[15] ), .Y(
        OR4_2596_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[20]  (.A(CFG3_12_Y), .B(
        CFG3_21_Y), .Y(\BLKY2[20] ));
    OR4 OR4_2797 (.A(\A_DOUT_TEMPR95[15] ), .B(\A_DOUT_TEMPR96[15] ), 
        .C(\A_DOUT_TEMPR97[15] ), .D(\A_DOUT_TEMPR98[15] ), .Y(
        OR4_2797_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%103%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R103C6 (
        .A_DOUT({nc27330, nc27331, nc27332, nc27333, nc27334, nc27335, 
        nc27336, nc27337, nc27338, nc27339, nc27340, nc27341, nc27342, 
        nc27343, nc27344, \A_DOUT_TEMPR103[34] , \A_DOUT_TEMPR103[33] , 
        \A_DOUT_TEMPR103[32] , \A_DOUT_TEMPR103[31] , 
        \A_DOUT_TEMPR103[30] }), .B_DOUT({nc27345, nc27346, nc27347, 
        nc27348, nc27349, nc27350, nc27351, nc27352, nc27353, nc27354, 
        nc27355, nc27356, nc27357, nc27358, nc27359, 
        \B_DOUT_TEMPR103[34] , \B_DOUT_TEMPR103[33] , 
        \B_DOUT_TEMPR103[32] , \B_DOUT_TEMPR103[31] , 
        \B_DOUT_TEMPR103[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[103][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2591 (.A(\A_DOUT_TEMPR0[39] ), .B(\A_DOUT_TEMPR1[39] ), .C(
        \A_DOUT_TEMPR2[39] ), .D(\A_DOUT_TEMPR3[39] ), .Y(OR4_2591_Y));
    OR4 OR4_955 (.A(\B_DOUT_TEMPR64[17] ), .B(\B_DOUT_TEMPR65[17] ), 
        .C(\B_DOUT_TEMPR66[17] ), .D(\B_DOUT_TEMPR67[17] ), .Y(
        OR4_955_Y));
    OR4 OR4_2770 (.A(OR4_1150_Y), .B(OR4_885_Y), .C(OR4_914_Y), .D(
        OR4_478_Y), .Y(OR4_2770_Y));
    OR4 OR4_455 (.A(\A_DOUT_TEMPR83[5] ), .B(\A_DOUT_TEMPR84[5] ), .C(
        \A_DOUT_TEMPR85[5] ), .D(\A_DOUT_TEMPR86[5] ), .Y(OR4_455_Y));
    OR4 OR4_1305 (.A(\A_DOUT_TEMPR60[35] ), .B(\A_DOUT_TEMPR61[35] ), 
        .C(\A_DOUT_TEMPR62[35] ), .D(\A_DOUT_TEMPR63[35] ), .Y(
        OR4_1305_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%21%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R21C2 (
        .A_DOUT({nc27360, nc27361, nc27362, nc27363, nc27364, nc27365, 
        nc27366, nc27367, nc27368, nc27369, nc27370, nc27371, nc27372, 
        nc27373, nc27374, \A_DOUT_TEMPR21[14] , \A_DOUT_TEMPR21[13] , 
        \A_DOUT_TEMPR21[12] , \A_DOUT_TEMPR21[11] , 
        \A_DOUT_TEMPR21[10] }), .B_DOUT({nc27375, nc27376, nc27377, 
        nc27378, nc27379, nc27380, nc27381, nc27382, nc27383, nc27384, 
        nc27385, nc27386, nc27387, nc27388, nc27389, 
        \B_DOUT_TEMPR21[14] , \B_DOUT_TEMPR21[13] , 
        \B_DOUT_TEMPR21[12] , \B_DOUT_TEMPR21[11] , 
        \B_DOUT_TEMPR21[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[21][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2351 (.A(OR4_2908_Y), .B(OR4_2625_Y), .C(OR4_1084_Y), .D(
        OR4_2631_Y), .Y(OR4_2351_Y));
    OR4 OR4_110 (.A(\B_DOUT_TEMPR24[11] ), .B(\B_DOUT_TEMPR25[11] ), 
        .C(\B_DOUT_TEMPR26[11] ), .D(\B_DOUT_TEMPR27[11] ), .Y(
        OR4_110_Y));
    OR4 OR4_887 (.A(\B_DOUT_TEMPR40[18] ), .B(\B_DOUT_TEMPR41[18] ), 
        .C(\B_DOUT_TEMPR42[18] ), .D(\B_DOUT_TEMPR43[18] ), .Y(
        OR4_887_Y));
    OR4 OR4_2851 (.A(\A_DOUT_TEMPR0[21] ), .B(\A_DOUT_TEMPR1[21] ), .C(
        \A_DOUT_TEMPR2[21] ), .D(\A_DOUT_TEMPR3[21] ), .Y(OR4_2851_Y));
    OR4 OR4_2586 (.A(OR4_1709_Y), .B(OR4_2538_Y), .C(OR2_39_Y), .D(
        \A_DOUT_TEMPR74[21] ), .Y(OR4_2586_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%80%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R80C7 (
        .A_DOUT({nc27390, nc27391, nc27392, nc27393, nc27394, nc27395, 
        nc27396, nc27397, nc27398, nc27399, nc27400, nc27401, nc27402, 
        nc27403, nc27404, \A_DOUT_TEMPR80[39] , \A_DOUT_TEMPR80[38] , 
        \A_DOUT_TEMPR80[37] , \A_DOUT_TEMPR80[36] , 
        \A_DOUT_TEMPR80[35] }), .B_DOUT({nc27405, nc27406, nc27407, 
        nc27408, nc27409, nc27410, nc27411, nc27412, nc27413, nc27414, 
        nc27415, nc27416, nc27417, nc27418, nc27419, 
        \B_DOUT_TEMPR80[39] , \B_DOUT_TEMPR80[38] , 
        \B_DOUT_TEMPR80[37] , \B_DOUT_TEMPR80[36] , 
        \B_DOUT_TEMPR80[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[80][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2440 (.A(\B_DOUT_TEMPR20[7] ), .B(\B_DOUT_TEMPR21[7] ), .C(
        \B_DOUT_TEMPR22[7] ), .D(\B_DOUT_TEMPR23[7] ), .Y(OR4_2440_Y));
    OR4 OR4_1750 (.A(\A_DOUT_TEMPR0[33] ), .B(\A_DOUT_TEMPR1[33] ), .C(
        \A_DOUT_TEMPR2[33] ), .D(\A_DOUT_TEMPR3[33] ), .Y(OR4_1750_Y));
    OR4 OR4_2787 (.A(\A_DOUT_TEMPR56[25] ), .B(\A_DOUT_TEMPR57[25] ), 
        .C(\A_DOUT_TEMPR58[25] ), .D(\A_DOUT_TEMPR59[25] ), .Y(
        OR4_2787_Y));
    OR4 OR4_2109 (.A(\A_DOUT_TEMPR48[38] ), .B(\A_DOUT_TEMPR49[38] ), 
        .C(\A_DOUT_TEMPR50[38] ), .D(\A_DOUT_TEMPR51[38] ), .Y(
        OR4_2109_Y));
    OR4 OR4_90 (.A(\A_DOUT_TEMPR103[12] ), .B(\A_DOUT_TEMPR104[12] ), 
        .C(\A_DOUT_TEMPR105[12] ), .D(\A_DOUT_TEMPR106[12] ), .Y(
        OR4_90_Y));
    OR4 OR4_2581 (.A(\B_DOUT_TEMPR115[9] ), .B(\B_DOUT_TEMPR116[9] ), 
        .C(\B_DOUT_TEMPR117[9] ), .D(\B_DOUT_TEMPR118[9] ), .Y(
        OR4_2581_Y));
    OR4 OR4_2466 (.A(OR4_2039_Y), .B(OR4_1273_Y), .C(OR4_1038_Y), .D(
        OR4_522_Y), .Y(OR4_2466_Y));
    CFG3 #( .INIT(8'h1) )  CFG3_11 (.A(B_ADDR[16]), .B(B_ADDR[15]), .C(
        B_ADDR[14]), .Y(CFG3_11_Y));
    OR4 OR4_618 (.A(\A_DOUT_TEMPR8[25] ), .B(\A_DOUT_TEMPR9[25] ), .C(
        \A_DOUT_TEMPR10[25] ), .D(\A_DOUT_TEMPR11[25] ), .Y(OR4_618_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%96%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R96C3 (
        .A_DOUT({nc27420, nc27421, nc27422, nc27423, nc27424, nc27425, 
        nc27426, nc27427, nc27428, nc27429, nc27430, nc27431, nc27432, 
        nc27433, nc27434, \A_DOUT_TEMPR96[19] , \A_DOUT_TEMPR96[18] , 
        \A_DOUT_TEMPR96[17] , \A_DOUT_TEMPR96[16] , 
        \A_DOUT_TEMPR96[15] }), .B_DOUT({nc27435, nc27436, nc27437, 
        nc27438, nc27439, nc27440, nc27441, nc27442, nc27443, nc27444, 
        nc27445, nc27446, nc27447, nc27448, nc27449, 
        \B_DOUT_TEMPR96[19] , \B_DOUT_TEMPR96[18] , 
        \B_DOUT_TEMPR96[17] , \B_DOUT_TEMPR96[16] , 
        \B_DOUT_TEMPR96[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[96][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2537 (.A(OR4_1400_Y), .B(OR4_1684_Y), .C(OR4_1348_Y), .D(
        OR4_1700_Y), .Y(OR4_2537_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%51%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R51C5 (
        .A_DOUT({nc27450, nc27451, nc27452, nc27453, nc27454, nc27455, 
        nc27456, nc27457, nc27458, nc27459, nc27460, nc27461, nc27462, 
        nc27463, nc27464, \A_DOUT_TEMPR51[29] , \A_DOUT_TEMPR51[28] , 
        \A_DOUT_TEMPR51[27] , \A_DOUT_TEMPR51[26] , 
        \A_DOUT_TEMPR51[25] }), .B_DOUT({nc27465, nc27466, nc27467, 
        nc27468, nc27469, nc27470, nc27471, nc27472, nc27473, nc27474, 
        nc27475, nc27476, nc27477, nc27478, nc27479, 
        \B_DOUT_TEMPR51[29] , \B_DOUT_TEMPR51[28] , 
        \B_DOUT_TEMPR51[27] , \B_DOUT_TEMPR51[26] , 
        \B_DOUT_TEMPR51[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[51][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[12] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[12] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2377 (.A(\B_DOUT_TEMPR40[31] ), .B(\B_DOUT_TEMPR41[31] ), 
        .C(\B_DOUT_TEMPR42[31] ), .D(\B_DOUT_TEMPR43[31] ), .Y(
        OR4_2377_Y));
    OR4 OR4_2272 (.A(OR4_2154_Y), .B(OR4_699_Y), .C(OR4_1523_Y), .D(
        OR4_552_Y), .Y(OR4_2272_Y));
    OR4 OR4_679 (.A(\B_DOUT_TEMPR115[3] ), .B(\B_DOUT_TEMPR116[3] ), 
        .C(\B_DOUT_TEMPR117[3] ), .D(\B_DOUT_TEMPR118[3] ), .Y(
        OR4_679_Y));
    OR4 OR4_1537 (.A(\B_DOUT_TEMPR48[29] ), .B(\B_DOUT_TEMPR49[29] ), 
        .C(\B_DOUT_TEMPR50[29] ), .D(\B_DOUT_TEMPR51[29] ), .Y(
        OR4_1537_Y));
    OR4 OR4_2245 (.A(\A_DOUT_TEMPR99[12] ), .B(\A_DOUT_TEMPR100[12] ), 
        .C(\A_DOUT_TEMPR101[12] ), .D(\A_DOUT_TEMPR102[12] ), .Y(
        OR4_2245_Y));
    OR4 OR4_1889 (.A(\B_DOUT_TEMPR99[8] ), .B(\B_DOUT_TEMPR100[8] ), 
        .C(\B_DOUT_TEMPR101[8] ), .D(\B_DOUT_TEMPR102[8] ), .Y(
        OR4_1889_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%47%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R47C4 (
        .A_DOUT({nc27480, nc27481, nc27482, nc27483, nc27484, nc27485, 
        nc27486, nc27487, nc27488, nc27489, nc27490, nc27491, nc27492, 
        nc27493, nc27494, \A_DOUT_TEMPR47[24] , \A_DOUT_TEMPR47[23] , 
        \A_DOUT_TEMPR47[22] , \A_DOUT_TEMPR47[21] , 
        \A_DOUT_TEMPR47[20] }), .B_DOUT({nc27495, nc27496, nc27497, 
        nc27498, nc27499, nc27500, nc27501, nc27502, nc27503, nc27504, 
        nc27505, nc27506, nc27507, nc27508, nc27509, 
        \B_DOUT_TEMPR47[24] , \B_DOUT_TEMPR47[23] , 
        \B_DOUT_TEMPR47[22] , \B_DOUT_TEMPR47[21] , 
        \B_DOUT_TEMPR47[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[47][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1943 (.A(\B_DOUT_TEMPR64[0] ), .B(\B_DOUT_TEMPR65[0] ), .C(
        \B_DOUT_TEMPR66[0] ), .D(\B_DOUT_TEMPR67[0] ), .Y(OR4_1943_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%5%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R5C3 (
        .A_DOUT({nc27510, nc27511, nc27512, nc27513, nc27514, nc27515, 
        nc27516, nc27517, nc27518, nc27519, nc27520, nc27521, nc27522, 
        nc27523, nc27524, \A_DOUT_TEMPR5[19] , \A_DOUT_TEMPR5[18] , 
        \A_DOUT_TEMPR5[17] , \A_DOUT_TEMPR5[16] , \A_DOUT_TEMPR5[15] })
        , .B_DOUT({nc27525, nc27526, nc27527, nc27528, nc27529, 
        nc27530, nc27531, nc27532, nc27533, nc27534, nc27535, nc27536, 
        nc27537, nc27538, nc27539, \B_DOUT_TEMPR5[19] , 
        \B_DOUT_TEMPR5[18] , \B_DOUT_TEMPR5[17] , \B_DOUT_TEMPR5[16] , 
        \B_DOUT_TEMPR5[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[5][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[1] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1665 (.A(\A_DOUT_TEMPR12[34] ), .B(\A_DOUT_TEMPR13[34] ), 
        .C(\A_DOUT_TEMPR14[34] ), .D(\A_DOUT_TEMPR15[34] ), .Y(
        OR4_1665_Y));
    OR4 OR4_2765 (.A(\A_DOUT_TEMPR44[36] ), .B(\A_DOUT_TEMPR45[36] ), 
        .C(\A_DOUT_TEMPR46[36] ), .D(\A_DOUT_TEMPR47[36] ), .Y(
        OR4_2765_Y));
    OR4 \OR4_B_DOUT[23]  (.A(OR4_829_Y), .B(OR4_543_Y), .C(OR4_2683_Y), 
        .D(OR4_232_Y), .Y(B_DOUT[23]));
    OR4 OR4_946 (.A(\A_DOUT_TEMPR44[5] ), .B(\A_DOUT_TEMPR45[5] ), .C(
        \A_DOUT_TEMPR46[5] ), .D(\A_DOUT_TEMPR47[5] ), .Y(OR4_946_Y));
    OR4 OR4_893 (.A(\A_DOUT_TEMPR99[7] ), .B(\A_DOUT_TEMPR100[7] ), .C(
        \A_DOUT_TEMPR101[7] ), .D(\A_DOUT_TEMPR102[7] ), .Y(OR4_893_Y));
    OR4 OR4_911 (.A(\A_DOUT_TEMPR52[17] ), .B(\A_DOUT_TEMPR53[17] ), 
        .C(\A_DOUT_TEMPR54[17] ), .D(\A_DOUT_TEMPR55[17] ), .Y(
        OR4_911_Y));
    OR4 OR4_1576 (.A(\A_DOUT_TEMPR0[13] ), .B(\A_DOUT_TEMPR1[13] ), .C(
        \A_DOUT_TEMPR2[13] ), .D(\A_DOUT_TEMPR3[13] ), .Y(OR4_1576_Y));
    OR4 OR4_1181 (.A(\B_DOUT_TEMPR16[6] ), .B(\B_DOUT_TEMPR17[6] ), .C(
        \B_DOUT_TEMPR18[6] ), .D(\B_DOUT_TEMPR19[6] ), .Y(OR4_1181_Y));
    OR4 OR4_1097 (.A(\A_DOUT_TEMPR68[9] ), .B(\A_DOUT_TEMPR69[9] ), .C(
        \A_DOUT_TEMPR70[9] ), .D(\A_DOUT_TEMPR71[9] ), .Y(OR4_1097_Y));
    OR4 OR4_1357 (.A(OR4_2672_Y), .B(OR4_810_Y), .C(OR2_45_Y), .D(
        \A_DOUT_TEMPR74[12] ), .Y(OR4_1357_Y));
    OR4 OR4_973 (.A(\A_DOUT_TEMPR4[36] ), .B(\A_DOUT_TEMPR5[36] ), .C(
        \A_DOUT_TEMPR6[36] ), .D(\A_DOUT_TEMPR7[36] ), .Y(OR4_973_Y));
    OR4 OR4_1252 (.A(\B_DOUT_TEMPR68[9] ), .B(\B_DOUT_TEMPR69[9] ), .C(
        \B_DOUT_TEMPR70[9] ), .D(\B_DOUT_TEMPR71[9] ), .Y(OR4_1252_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%22%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R22C3 (
        .A_DOUT({nc27540, nc27541, nc27542, nc27543, nc27544, nc27545, 
        nc27546, nc27547, nc27548, nc27549, nc27550, nc27551, nc27552, 
        nc27553, nc27554, \A_DOUT_TEMPR22[19] , \A_DOUT_TEMPR22[18] , 
        \A_DOUT_TEMPR22[17] , \A_DOUT_TEMPR22[16] , 
        \A_DOUT_TEMPR22[15] }), .B_DOUT({nc27555, nc27556, nc27557, 
        nc27558, nc27559, nc27560, nc27561, nc27562, nc27563, nc27564, 
        nc27565, nc27566, nc27567, nc27568, nc27569, 
        \B_DOUT_TEMPR22[19] , \B_DOUT_TEMPR22[18] , 
        \B_DOUT_TEMPR22[17] , \B_DOUT_TEMPR22[16] , 
        \B_DOUT_TEMPR22[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[22][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1399 (.A(\B_DOUT_TEMPR115[25] ), .B(\B_DOUT_TEMPR116[25] ), 
        .C(\B_DOUT_TEMPR117[25] ), .D(\B_DOUT_TEMPR118[25] ), .Y(
        OR4_1399_Y));
    OR4 OR4_1777 (.A(\B_DOUT_TEMPR99[15] ), .B(\B_DOUT_TEMPR100[15] ), 
        .C(\B_DOUT_TEMPR101[15] ), .D(\B_DOUT_TEMPR102[15] ), .Y(
        OR4_1777_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%43%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R43C6 (
        .A_DOUT({nc27570, nc27571, nc27572, nc27573, nc27574, nc27575, 
        nc27576, nc27577, nc27578, nc27579, nc27580, nc27581, nc27582, 
        nc27583, nc27584, \A_DOUT_TEMPR43[34] , \A_DOUT_TEMPR43[33] , 
        \A_DOUT_TEMPR43[32] , \A_DOUT_TEMPR43[31] , 
        \A_DOUT_TEMPR43[30] }), .B_DOUT({nc27585, nc27586, nc27587, 
        nc27588, nc27589, nc27590, nc27591, nc27592, nc27593, nc27594, 
        nc27595, nc27596, nc27597, nc27598, nc27599, 
        \B_DOUT_TEMPR43[34] , \B_DOUT_TEMPR43[33] , 
        \B_DOUT_TEMPR43[32] , \B_DOUT_TEMPR43[31] , 
        \B_DOUT_TEMPR43[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[43][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2474 (.A(\B_DOUT_TEMPR16[11] ), .B(\B_DOUT_TEMPR17[11] ), 
        .C(\B_DOUT_TEMPR18[11] ), .D(\B_DOUT_TEMPR19[11] ), .Y(
        OR4_2474_Y));
    OR4 OR4_1341 (.A(\A_DOUT_TEMPR16[34] ), .B(\A_DOUT_TEMPR17[34] ), 
        .C(\A_DOUT_TEMPR18[34] ), .D(\A_DOUT_TEMPR19[34] ), .Y(
        OR4_1341_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%20%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R20C3 (
        .A_DOUT({nc27600, nc27601, nc27602, nc27603, nc27604, nc27605, 
        nc27606, nc27607, nc27608, nc27609, nc27610, nc27611, nc27612, 
        nc27613, nc27614, \A_DOUT_TEMPR20[19] , \A_DOUT_TEMPR20[18] , 
        \A_DOUT_TEMPR20[17] , \A_DOUT_TEMPR20[16] , 
        \A_DOUT_TEMPR20[15] }), .B_DOUT({nc27615, nc27616, nc27617, 
        nc27618, nc27619, nc27620, nc27621, nc27622, nc27623, nc27624, 
        nc27625, nc27626, nc27627, nc27628, nc27629, 
        \B_DOUT_TEMPR20[19] , \B_DOUT_TEMPR20[18] , 
        \B_DOUT_TEMPR20[17] , \B_DOUT_TEMPR20[16] , 
        \B_DOUT_TEMPR20[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[20][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1297 (.A(\A_DOUT_TEMPR75[31] ), .B(\A_DOUT_TEMPR76[31] ), 
        .C(\A_DOUT_TEMPR77[31] ), .D(\A_DOUT_TEMPR78[31] ), .Y(
        OR4_1297_Y));
    OR4 OR4_1571 (.A(OR4_1701_Y), .B(OR4_1076_Y), .C(OR4_575_Y), .D(
        OR4_882_Y), .Y(OR4_1571_Y));
    OR4 OR4_1085 (.A(\A_DOUT_TEMPR115[33] ), .B(\A_DOUT_TEMPR116[33] ), 
        .C(\A_DOUT_TEMPR117[33] ), .D(\A_DOUT_TEMPR118[33] ), .Y(
        OR4_1085_Y));
    OR4 OR4_1667 (.A(\A_DOUT_TEMPR99[27] ), .B(\A_DOUT_TEMPR100[27] ), 
        .C(\A_DOUT_TEMPR101[27] ), .D(\A_DOUT_TEMPR102[27] ), .Y(
        OR4_1667_Y));
    OR4 OR4_1841 (.A(OR4_648_Y), .B(OR4_447_Y), .C(OR4_1336_Y), .D(
        OR4_2509_Y), .Y(OR4_1841_Y));
    OR4 OR4_422 (.A(\B_DOUT_TEMPR36[32] ), .B(\B_DOUT_TEMPR37[32] ), 
        .C(\B_DOUT_TEMPR38[32] ), .D(\B_DOUT_TEMPR39[32] ), .Y(
        OR4_422_Y));
    OR4 OR4_1990 (.A(\B_DOUT_TEMPR48[8] ), .B(\B_DOUT_TEMPR49[8] ), .C(
        \B_DOUT_TEMPR50[8] ), .D(\B_DOUT_TEMPR51[8] ), .Y(OR4_1990_Y));
    OR4 OR4_192 (.A(\A_DOUT_TEMPR111[31] ), .B(\A_DOUT_TEMPR112[31] ), 
        .C(\A_DOUT_TEMPR113[31] ), .D(\A_DOUT_TEMPR114[31] ), .Y(
        OR4_192_Y));
    OR4 OR4_1220 (.A(OR4_738_Y), .B(OR4_1116_Y), .C(OR4_1719_Y), .D(
        OR4_950_Y), .Y(OR4_1220_Y));
    OR4 OR4_2829 (.A(\A_DOUT_TEMPR107[28] ), .B(\A_DOUT_TEMPR108[28] ), 
        .C(\A_DOUT_TEMPR109[28] ), .D(\A_DOUT_TEMPR110[28] ), .Y(
        OR4_2829_Y));
    OR4 OR4_77 (.A(OR4_2954_Y), .B(OR4_33_Y), .C(OR4_657_Y), .D(
        OR4_2902_Y), .Y(OR4_77_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%109%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R109C7 (
        .A_DOUT({nc27630, nc27631, nc27632, nc27633, nc27634, nc27635, 
        nc27636, nc27637, nc27638, nc27639, nc27640, nc27641, nc27642, 
        nc27643, nc27644, \A_DOUT_TEMPR109[39] , \A_DOUT_TEMPR109[38] , 
        \A_DOUT_TEMPR109[37] , \A_DOUT_TEMPR109[36] , 
        \A_DOUT_TEMPR109[35] }), .B_DOUT({nc27645, nc27646, nc27647, 
        nc27648, nc27649, nc27650, nc27651, nc27652, nc27653, nc27654, 
        nc27655, nc27656, nc27657, nc27658, nc27659, 
        \B_DOUT_TEMPR109[39] , \B_DOUT_TEMPR109[38] , 
        \B_DOUT_TEMPR109[37] , \B_DOUT_TEMPR109[36] , 
        \B_DOUT_TEMPR109[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[109][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%26%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R26C6 (
        .A_DOUT({nc27660, nc27661, nc27662, nc27663, nc27664, nc27665, 
        nc27666, nc27667, nc27668, nc27669, nc27670, nc27671, nc27672, 
        nc27673, nc27674, \A_DOUT_TEMPR26[34] , \A_DOUT_TEMPR26[33] , 
        \A_DOUT_TEMPR26[32] , \A_DOUT_TEMPR26[31] , 
        \A_DOUT_TEMPR26[30] }), .B_DOUT({nc27675, nc27676, nc27677, 
        nc27678, nc27679, nc27680, nc27681, nc27682, nc27683, nc27684, 
        nc27685, nc27686, nc27687, nc27688, nc27689, 
        \B_DOUT_TEMPR26[34] , \B_DOUT_TEMPR26[33] , 
        \B_DOUT_TEMPR26[32] , \B_DOUT_TEMPR26[31] , 
        \B_DOUT_TEMPR26[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], B_DIN[32], 
        B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1454 (.A(\B_DOUT_TEMPR40[3] ), .B(\B_DOUT_TEMPR41[3] ), .C(
        \B_DOUT_TEMPR42[3] ), .D(\B_DOUT_TEMPR43[3] ), .Y(OR4_1454_Y));
    OR4 OR4_609 (.A(OR4_2387_Y), .B(OR4_1419_Y), .C(OR4_1618_Y), .D(
        OR4_1428_Y), .Y(OR4_609_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%71%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R71C0 (
        .A_DOUT({nc27690, nc27691, nc27692, nc27693, nc27694, nc27695, 
        nc27696, nc27697, nc27698, nc27699, nc27700, nc27701, nc27702, 
        nc27703, nc27704, \A_DOUT_TEMPR71[4] , \A_DOUT_TEMPR71[3] , 
        \A_DOUT_TEMPR71[2] , \A_DOUT_TEMPR71[1] , \A_DOUT_TEMPR71[0] })
        , .B_DOUT({nc27705, nc27706, nc27707, nc27708, nc27709, 
        nc27710, nc27711, nc27712, nc27713, nc27714, nc27715, nc27716, 
        nc27717, nc27718, nc27719, \B_DOUT_TEMPR71[4] , 
        \B_DOUT_TEMPR71[3] , \B_DOUT_TEMPR71[2] , \B_DOUT_TEMPR71[1] , 
        \B_DOUT_TEMPR71[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[71][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[17] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[17] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_481 (.A(\B_DOUT_TEMPR79[30] ), .B(\B_DOUT_TEMPR80[30] ), 
        .C(\B_DOUT_TEMPR81[30] ), .D(\B_DOUT_TEMPR82[30] ), .Y(
        OR4_481_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%82%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R82C0 (
        .A_DOUT({nc27720, nc27721, nc27722, nc27723, nc27724, nc27725, 
        nc27726, nc27727, nc27728, nc27729, nc27730, nc27731, nc27732, 
        nc27733, nc27734, \A_DOUT_TEMPR82[4] , \A_DOUT_TEMPR82[3] , 
        \A_DOUT_TEMPR82[2] , \A_DOUT_TEMPR82[1] , \A_DOUT_TEMPR82[0] })
        , .B_DOUT({nc27735, nc27736, nc27737, nc27738, nc27739, 
        nc27740, nc27741, nc27742, nc27743, nc27744, nc27745, nc27746, 
        nc27747, nc27748, nc27749, \B_DOUT_TEMPR82[4] , 
        \B_DOUT_TEMPR82[3] , \B_DOUT_TEMPR82[2] , \B_DOUT_TEMPR82[1] , 
        \B_DOUT_TEMPR82[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[82][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%31%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R31C5 (
        .A_DOUT({nc27750, nc27751, nc27752, nc27753, nc27754, nc27755, 
        nc27756, nc27757, nc27758, nc27759, nc27760, nc27761, nc27762, 
        nc27763, nc27764, \A_DOUT_TEMPR31[29] , \A_DOUT_TEMPR31[28] , 
        \A_DOUT_TEMPR31[27] , \A_DOUT_TEMPR31[26] , 
        \A_DOUT_TEMPR31[25] }), .B_DOUT({nc27765, nc27766, nc27767, 
        nc27768, nc27769, nc27770, nc27771, nc27772, nc27773, nc27774, 
        nc27775, nc27776, nc27777, nc27778, nc27779, 
        \B_DOUT_TEMPR31[29] , \B_DOUT_TEMPR31[28] , 
        \B_DOUT_TEMPR31[27] , \B_DOUT_TEMPR31[26] , 
        \B_DOUT_TEMPR31[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[31][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[7] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[7] , B_ADDR[13], B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], B_DIN[27], 
        B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1917 (.A(\B_DOUT_TEMPR95[10] ), .B(\B_DOUT_TEMPR96[10] ), 
        .C(\B_DOUT_TEMPR97[10] ), .D(\B_DOUT_TEMPR98[10] ), .Y(
        OR4_1917_Y));
    OR4 OR4_1887 (.A(\B_DOUT_TEMPR95[4] ), .B(\B_DOUT_TEMPR96[4] ), .C(
        \B_DOUT_TEMPR97[4] ), .D(\B_DOUT_TEMPR98[4] ), .Y(OR4_1887_Y));
    OR4 OR4_2238 (.A(\A_DOUT_TEMPR12[1] ), .B(\A_DOUT_TEMPR13[1] ), .C(
        \A_DOUT_TEMPR14[1] ), .D(\A_DOUT_TEMPR15[1] ), .Y(OR4_2238_Y));
    OR4 OR4_914 (.A(OR4_706_Y), .B(OR4_1639_Y), .C(OR4_2271_Y), .D(
        OR4_1463_Y), .Y(OR4_914_Y));
    OR4 OR4_995 (.A(\B_DOUT_TEMPR99[9] ), .B(\B_DOUT_TEMPR100[9] ), .C(
        \B_DOUT_TEMPR101[9] ), .D(\B_DOUT_TEMPR102[9] ), .Y(OR4_995_Y));
    OR4 OR4_495 (.A(\A_DOUT_TEMPR115[30] ), .B(\A_DOUT_TEMPR116[30] ), 
        .C(\A_DOUT_TEMPR117[30] ), .D(\A_DOUT_TEMPR118[30] ), .Y(
        OR4_495_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[24]  (.A(CFG3_17_Y), .B(
        CFG3_18_Y), .Y(\BLKX2[24] ));
    OR4 OR4_2121 (.A(\A_DOUT_TEMPR8[9] ), .B(\A_DOUT_TEMPR9[9] ), .C(
        \A_DOUT_TEMPR10[9] ), .D(\A_DOUT_TEMPR11[9] ), .Y(OR4_2121_Y));
    OR4 OR4_1238 (.A(\B_DOUT_TEMPR8[0] ), .B(\B_DOUT_TEMPR9[0] ), .C(
        \B_DOUT_TEMPR10[0] ), .D(\B_DOUT_TEMPR11[0] ), .Y(OR4_1238_Y));
    OR4 OR4_1792 (.A(\A_DOUT_TEMPR40[22] ), .B(\A_DOUT_TEMPR41[22] ), 
        .C(\A_DOUT_TEMPR42[22] ), .D(\A_DOUT_TEMPR43[22] ), .Y(
        OR4_1792_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%107%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R107C1 (
        .A_DOUT({nc27780, nc27781, nc27782, nc27783, nc27784, nc27785, 
        nc27786, nc27787, nc27788, nc27789, nc27790, nc27791, nc27792, 
        nc27793, nc27794, \A_DOUT_TEMPR107[9] , \A_DOUT_TEMPR107[8] , 
        \A_DOUT_TEMPR107[7] , \A_DOUT_TEMPR107[6] , 
        \A_DOUT_TEMPR107[5] }), .B_DOUT({nc27795, nc27796, nc27797, 
        nc27798, nc27799, nc27800, nc27801, nc27802, nc27803, nc27804, 
        nc27805, nc27806, nc27807, nc27808, nc27809, 
        \B_DOUT_TEMPR107[9] , \B_DOUT_TEMPR107[8] , 
        \B_DOUT_TEMPR107[7] , \B_DOUT_TEMPR107[6] , 
        \B_DOUT_TEMPR107[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[107][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%81%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R81C6 (
        .A_DOUT({nc27810, nc27811, nc27812, nc27813, nc27814, nc27815, 
        nc27816, nc27817, nc27818, nc27819, nc27820, nc27821, nc27822, 
        nc27823, nc27824, \A_DOUT_TEMPR81[34] , \A_DOUT_TEMPR81[33] , 
        \A_DOUT_TEMPR81[32] , \A_DOUT_TEMPR81[31] , 
        \A_DOUT_TEMPR81[30] }), .B_DOUT({nc27825, nc27826, nc27827, 
        nc27828, nc27829, nc27830, nc27831, nc27832, nc27833, nc27834, 
        nc27835, nc27836, nc27837, nc27838, nc27839, 
        \B_DOUT_TEMPR81[34] , \B_DOUT_TEMPR81[33] , 
        \B_DOUT_TEMPR81[32] , \B_DOUT_TEMPR81[31] , 
        \B_DOUT_TEMPR81[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[81][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2898 (.A(OR4_1172_Y), .B(OR4_843_Y), .C(OR4_1462_Y), .D(
        OR4_663_Y), .Y(OR4_2898_Y));
    OR4 OR4_2802 (.A(\A_DOUT_TEMPR87[6] ), .B(\A_DOUT_TEMPR88[6] ), .C(
        \A_DOUT_TEMPR89[6] ), .D(\A_DOUT_TEMPR90[6] ), .Y(OR4_2802_Y));
    OR4 OR4_1326 (.A(\A_DOUT_TEMPR48[36] ), .B(\A_DOUT_TEMPR49[36] ), 
        .C(\A_DOUT_TEMPR50[36] ), .D(\A_DOUT_TEMPR51[36] ), .Y(
        OR4_1326_Y));
    OR4 OR4_903 (.A(OR4_2349_Y), .B(OR4_258_Y), .C(OR4_2443_Y), .D(
        OR4_2813_Y), .Y(OR4_903_Y));
    OR4 OR4_95 (.A(\A_DOUT_TEMPR20[14] ), .B(\A_DOUT_TEMPR21[14] ), .C(
        \A_DOUT_TEMPR22[14] ), .D(\A_DOUT_TEMPR23[14] ), .Y(OR4_95_Y));
    OR4 OR4_2025 (.A(OR4_607_Y), .B(OR4_2307_Y), .C(OR4_1213_Y), .D(
        OR4_1402_Y), .Y(OR4_2025_Y));
    OR4 OR4_2646 (.A(\A_DOUT_TEMPR99[1] ), .B(\A_DOUT_TEMPR100[1] ), 
        .C(\A_DOUT_TEMPR101[1] ), .D(\A_DOUT_TEMPR102[1] ), .Y(
        OR4_2646_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%114%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R114C2 (
        .A_DOUT({nc27840, nc27841, nc27842, nc27843, nc27844, nc27845, 
        nc27846, nc27847, nc27848, nc27849, nc27850, nc27851, nc27852, 
        nc27853, nc27854, \A_DOUT_TEMPR114[14] , \A_DOUT_TEMPR114[13] , 
        \A_DOUT_TEMPR114[12] , \A_DOUT_TEMPR114[11] , 
        \A_DOUT_TEMPR114[10] }), .B_DOUT({nc27855, nc27856, nc27857, 
        nc27858, nc27859, nc27860, nc27861, nc27862, nc27863, nc27864, 
        nc27865, nc27866, nc27867, nc27868, nc27869, 
        \B_DOUT_TEMPR114[14] , \B_DOUT_TEMPR114[13] , 
        \B_DOUT_TEMPR114[12] , \B_DOUT_TEMPR114[11] , 
        \B_DOUT_TEMPR114[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[114][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2140 (.A(OR4_2551_Y), .B(OR4_320_Y), .C(OR2_59_Y), .D(
        \A_DOUT_TEMPR74[24] ), .Y(OR4_2140_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%44%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R44C4 (
        .A_DOUT({nc27870, nc27871, nc27872, nc27873, nc27874, nc27875, 
        nc27876, nc27877, nc27878, nc27879, nc27880, nc27881, nc27882, 
        nc27883, nc27884, \A_DOUT_TEMPR44[24] , \A_DOUT_TEMPR44[23] , 
        \A_DOUT_TEMPR44[22] , \A_DOUT_TEMPR44[21] , 
        \A_DOUT_TEMPR44[20] }), .B_DOUT({nc27885, nc27886, nc27887, 
        nc27888, nc27889, nc27890, nc27891, nc27892, nc27893, nc27894, 
        nc27895, nc27896, nc27897, nc27898, nc27899, 
        \B_DOUT_TEMPR44[24] , \B_DOUT_TEMPR44[23] , 
        \B_DOUT_TEMPR44[22] , \B_DOUT_TEMPR44[21] , 
        \B_DOUT_TEMPR44[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[44][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%104%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R104C5 (
        .A_DOUT({nc27900, nc27901, nc27902, nc27903, nc27904, nc27905, 
        nc27906, nc27907, nc27908, nc27909, nc27910, nc27911, nc27912, 
        nc27913, nc27914, \A_DOUT_TEMPR104[29] , \A_DOUT_TEMPR104[28] , 
        \A_DOUT_TEMPR104[27] , \A_DOUT_TEMPR104[26] , 
        \A_DOUT_TEMPR104[25] }), .B_DOUT({nc27915, nc27916, nc27917, 
        nc27918, nc27919, nc27920, nc27921, nc27922, nc27923, nc27924, 
        nc27925, nc27926, nc27927, nc27928, nc27929, 
        \B_DOUT_TEMPR104[29] , \B_DOUT_TEMPR104[28] , 
        \B_DOUT_TEMPR104[27] , \B_DOUT_TEMPR104[26] , 
        \B_DOUT_TEMPR104[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[104][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1810 (.A(OR4_362_Y), .B(OR4_702_Y), .C(OR4_1401_Y), .D(
        OR4_1681_Y), .Y(OR4_1810_Y));
    OR4 OR4_160 (.A(OR4_107_Y), .B(OR4_2322_Y), .C(OR4_1328_Y), .D(
        OR4_1608_Y), .Y(OR4_160_Y));
    OR4 OR4_1 (.A(OR4_684_Y), .B(OR4_23_Y), .C(OR2_47_Y), .D(
        \B_DOUT_TEMPR74[4] ), .Y(OR4_1_Y));
    OR4 OR4_2274 (.A(\B_DOUT_TEMPR0[33] ), .B(\B_DOUT_TEMPR1[33] ), .C(
        \B_DOUT_TEMPR2[33] ), .D(\B_DOUT_TEMPR3[33] ), .Y(OR4_2274_Y));
    OR4 OR4_2957 (.A(\A_DOUT_TEMPR87[5] ), .B(\A_DOUT_TEMPR88[5] ), .C(
        \A_DOUT_TEMPR89[5] ), .D(\A_DOUT_TEMPR90[5] ), .Y(OR4_2957_Y));
    OR4 OR4_1692 (.A(\B_DOUT_TEMPR16[28] ), .B(\B_DOUT_TEMPR17[28] ), 
        .C(\B_DOUT_TEMPR18[28] ), .D(\B_DOUT_TEMPR19[28] ), .Y(
        OR4_1692_Y));
    OR4 OR4_1364 (.A(\A_DOUT_TEMPR12[31] ), .B(\A_DOUT_TEMPR13[31] ), 
        .C(\A_DOUT_TEMPR14[31] ), .D(\A_DOUT_TEMPR15[31] ), .Y(
        OR4_1364_Y));
    OR4 OR4_70 (.A(\B_DOUT_TEMPR20[32] ), .B(\B_DOUT_TEMPR21[32] ), .C(
        \B_DOUT_TEMPR22[32] ), .D(\B_DOUT_TEMPR23[32] ), .Y(OR4_70_Y));
    OR4 OR4_2888 (.A(OR4_2005_Y), .B(OR4_3003_Y), .C(OR4_637_Y), .D(
        OR4_2285_Y), .Y(OR4_2888_Y));
    OR4 OR4_2566 (.A(\B_DOUT_TEMPR56[12] ), .B(\B_DOUT_TEMPR57[12] ), 
        .C(\B_DOUT_TEMPR58[12] ), .D(\B_DOUT_TEMPR59[12] ), .Y(
        OR4_2566_Y));
    OR4 OR4_2827 (.A(\A_DOUT_TEMPR60[4] ), .B(\A_DOUT_TEMPR61[4] ), .C(
        \A_DOUT_TEMPR62[4] ), .D(\A_DOUT_TEMPR63[4] ), .Y(OR4_2827_Y));
    OR4 OR4_1814 (.A(\A_DOUT_TEMPR79[5] ), .B(\A_DOUT_TEMPR80[5] ), .C(
        \A_DOUT_TEMPR81[5] ), .D(\A_DOUT_TEMPR82[5] ), .Y(OR4_1814_Y));
    OR4 OR4_2603 (.A(\B_DOUT_TEMPR4[33] ), .B(\B_DOUT_TEMPR5[33] ), .C(
        \B_DOUT_TEMPR6[33] ), .D(\B_DOUT_TEMPR7[33] ), .Y(OR4_2603_Y));
    OR4 OR4_442 (.A(\A_DOUT_TEMPR83[26] ), .B(\A_DOUT_TEMPR84[26] ), 
        .C(\A_DOUT_TEMPR85[26] ), .D(\A_DOUT_TEMPR86[26] ), .Y(
        OR4_442_Y));
    OR4 OR4_2767 (.A(OR4_1022_Y), .B(OR4_2729_Y), .C(OR4_1164_Y), .D(
        OR4_2730_Y), .Y(OR4_2767_Y));
    OR4 OR4_1992 (.A(\A_DOUT_TEMPR8[29] ), .B(\A_DOUT_TEMPR9[29] ), .C(
        \A_DOUT_TEMPR10[29] ), .D(\A_DOUT_TEMPR11[29] ), .Y(OR4_1992_Y)
        );
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%90%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R90C0 (
        .A_DOUT({nc27930, nc27931, nc27932, nc27933, nc27934, nc27935, 
        nc27936, nc27937, nc27938, nc27939, nc27940, nc27941, nc27942, 
        nc27943, nc27944, \A_DOUT_TEMPR90[4] , \A_DOUT_TEMPR90[3] , 
        \A_DOUT_TEMPR90[2] , \A_DOUT_TEMPR90[1] , \A_DOUT_TEMPR90[0] })
        , .B_DOUT({nc27945, nc27946, nc27947, nc27948, nc27949, 
        nc27950, nc27951, nc27952, nc27953, nc27954, nc27955, nc27956, 
        nc27957, nc27958, nc27959, \B_DOUT_TEMPR90[4] , 
        \B_DOUT_TEMPR90[3] , \B_DOUT_TEMPR90[2] , \B_DOUT_TEMPR90[1] , 
        \B_DOUT_TEMPR90[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[90][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%9%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R9C2 (
        .A_DOUT({nc27960, nc27961, nc27962, nc27963, nc27964, nc27965, 
        nc27966, nc27967, nc27968, nc27969, nc27970, nc27971, nc27972, 
        nc27973, nc27974, \A_DOUT_TEMPR9[14] , \A_DOUT_TEMPR9[13] , 
        \A_DOUT_TEMPR9[12] , \A_DOUT_TEMPR9[11] , \A_DOUT_TEMPR9[10] })
        , .B_DOUT({nc27975, nc27976, nc27977, nc27978, nc27979, 
        nc27980, nc27981, nc27982, nc27983, nc27984, nc27985, nc27986, 
        nc27987, nc27988, nc27989, \B_DOUT_TEMPR9[14] , 
        \B_DOUT_TEMPR9[13] , \B_DOUT_TEMPR9[12] , \B_DOUT_TEMPR9[11] , 
        \B_DOUT_TEMPR9[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[9][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[2] , \BLKY1[0] , B_ADDR[12]}), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], B_DIN[12], 
        B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2909 (.A(OR4_371_Y), .B(OR4_1302_Y), .C(OR4_961_Y), .D(
        OR4_2424_Y), .Y(OR4_2909_Y));
    OR4 OR4_2561 (.A(\A_DOUT_TEMPR107[9] ), .B(\A_DOUT_TEMPR108[9] ), 
        .C(\A_DOUT_TEMPR109[9] ), .D(\A_DOUT_TEMPR110[9] ), .Y(
        OR4_2561_Y));
    OR4 OR4_668 (.A(\B_DOUT_TEMPR103[24] ), .B(\B_DOUT_TEMPR104[24] ), 
        .C(\B_DOUT_TEMPR105[24] ), .D(\B_DOUT_TEMPR106[24] ), .Y(
        OR4_668_Y));
    OR4 OR4_2073 (.A(\B_DOUT_TEMPR12[28] ), .B(\B_DOUT_TEMPR13[28] ), 
        .C(\B_DOUT_TEMPR14[28] ), .D(\B_DOUT_TEMPR15[28] ), .Y(
        OR4_2073_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%95%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R95C4 (
        .A_DOUT({nc27990, nc27991, nc27992, nc27993, nc27994, nc27995, 
        nc27996, nc27997, nc27998, nc27999, nc28000, nc28001, nc28002, 
        nc28003, nc28004, \A_DOUT_TEMPR95[24] , \A_DOUT_TEMPR95[23] , 
        \A_DOUT_TEMPR95[22] , \A_DOUT_TEMPR95[21] , 
        \A_DOUT_TEMPR95[20] }), .B_DOUT({nc28005, nc28006, nc28007, 
        nc28008, nc28009, nc28010, nc28011, nc28012, nc28013, nc28014, 
        nc28015, nc28016, nc28017, nc28018, nc28019, 
        \B_DOUT_TEMPR95[24] , \B_DOUT_TEMPR95[23] , 
        \B_DOUT_TEMPR95[22] , \B_DOUT_TEMPR95[21] , 
        \B_DOUT_TEMPR95[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[95][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[23] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[23] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1254 (.A(\A_DOUT_TEMPR91[16] ), .B(\A_DOUT_TEMPR92[16] ), 
        .C(\A_DOUT_TEMPR93[16] ), .D(\A_DOUT_TEMPR94[16] ), .Y(
        OR4_1254_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%107%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R107C0 (
        .A_DOUT({nc28020, nc28021, nc28022, nc28023, nc28024, nc28025, 
        nc28026, nc28027, nc28028, nc28029, nc28030, nc28031, nc28032, 
        nc28033, nc28034, \A_DOUT_TEMPR107[4] , \A_DOUT_TEMPR107[3] , 
        \A_DOUT_TEMPR107[2] , \A_DOUT_TEMPR107[1] , 
        \A_DOUT_TEMPR107[0] }), .B_DOUT({nc28035, nc28036, nc28037, 
        nc28038, nc28039, nc28040, nc28041, nc28042, nc28043, nc28044, 
        nc28045, nc28046, nc28047, nc28048, nc28049, 
        \B_DOUT_TEMPR107[4] , \B_DOUT_TEMPR107[3] , 
        \B_DOUT_TEMPR107[2] , \B_DOUT_TEMPR107[1] , 
        \B_DOUT_TEMPR107[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[107][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[26] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[26] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], 
        B_DIN[2], B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[0] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%88%2%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R88C2 (
        .A_DOUT({nc28050, nc28051, nc28052, nc28053, nc28054, nc28055, 
        nc28056, nc28057, nc28058, nc28059, nc28060, nc28061, nc28062, 
        nc28063, nc28064, \A_DOUT_TEMPR88[14] , \A_DOUT_TEMPR88[13] , 
        \A_DOUT_TEMPR88[12] , \A_DOUT_TEMPR88[11] , 
        \A_DOUT_TEMPR88[10] }), .B_DOUT({nc28065, nc28066, nc28067, 
        nc28068, nc28069, nc28070, nc28071, nc28072, nc28073, nc28074, 
        nc28075, nc28076, nc28077, nc28078, nc28079, 
        \B_DOUT_TEMPR88[14] , \B_DOUT_TEMPR88[13] , 
        \B_DOUT_TEMPR88[12] , \B_DOUT_TEMPR88[11] , 
        \B_DOUT_TEMPR88[10] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[88][2] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[14], 
        A_DIN[13], A_DIN[12], A_DIN[11], A_DIN[10]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[4] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[14], B_DIN[13], 
        B_DIN[12], B_DIN[11], B_DIN[10]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[4] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2671 (.A(OR4_1367_Y), .B(OR4_1641_Y), .C(OR4_1301_Y), .D(
        OR4_1662_Y), .Y(OR4_2671_Y));
    OR4 OR4_2850 (.A(OR4_1855_Y), .B(OR4_2687_Y), .C(OR2_43_Y), .D(
        \B_DOUT_TEMPR74[23] ), .Y(OR4_2850_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%110%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R110C7 (
        .A_DOUT({nc28080, nc28081, nc28082, nc28083, nc28084, nc28085, 
        nc28086, nc28087, nc28088, nc28089, nc28090, nc28091, nc28092, 
        nc28093, nc28094, \A_DOUT_TEMPR110[39] , \A_DOUT_TEMPR110[38] , 
        \A_DOUT_TEMPR110[37] , \A_DOUT_TEMPR110[36] , 
        \A_DOUT_TEMPR110[35] }), .B_DOUT({nc28095, nc28096, nc28097, 
        nc28098, nc28099, nc28100, nc28101, nc28102, nc28103, nc28104, 
        nc28105, nc28106, nc28107, nc28108, nc28109, 
        \B_DOUT_TEMPR110[39] , \B_DOUT_TEMPR110[38] , 
        \B_DOUT_TEMPR110[37] , \B_DOUT_TEMPR110[36] , 
        \B_DOUT_TEMPR110[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[110][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[27] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[27] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2773 (.A(OR4_517_Y), .B(OR4_2904_Y), .C(OR4_1756_Y), .D(
        OR4_1394_Y), .Y(OR4_2773_Y));
    OR4 OR4_2798 (.A(\B_DOUT_TEMPR83[12] ), .B(\B_DOUT_TEMPR84[12] ), 
        .C(\B_DOUT_TEMPR85[12] ), .D(\B_DOUT_TEMPR86[12] ), .Y(
        OR4_2798_Y));
    OR4 \OR4_A_DOUT[32]  (.A(OR4_661_Y), .B(OR4_2243_Y), .C(OR4_159_Y), 
        .D(OR4_2915_Y), .Y(A_DOUT[32]));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%56%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R56C3 (
        .A_DOUT({nc28110, nc28111, nc28112, nc28113, nc28114, nc28115, 
        nc28116, nc28117, nc28118, nc28119, nc28120, nc28121, nc28122, 
        nc28123, nc28124, \A_DOUT_TEMPR56[19] , \A_DOUT_TEMPR56[18] , 
        \A_DOUT_TEMPR56[17] , \A_DOUT_TEMPR56[16] , 
        \A_DOUT_TEMPR56[15] }), .B_DOUT({nc28125, nc28126, nc28127, 
        nc28128, nc28129, nc28130, nc28131, nc28132, nc28133, nc28134, 
        nc28135, nc28136, nc28137, nc28138, nc28139, 
        \B_DOUT_TEMPR56[19] , \B_DOUT_TEMPR56[18] , 
        \B_DOUT_TEMPR56[17] , \B_DOUT_TEMPR56[16] , 
        \B_DOUT_TEMPR56[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[56][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1503 (.A(\A_DOUT_TEMPR103[36] ), .B(\A_DOUT_TEMPR104[36] ), 
        .C(\A_DOUT_TEMPR105[36] ), .D(\A_DOUT_TEMPR106[36] ), .Y(
        OR4_1503_Y));
    OR4 OR4_2175 (.A(\A_DOUT_TEMPR60[13] ), .B(\A_DOUT_TEMPR61[13] ), 
        .C(\A_DOUT_TEMPR62[13] ), .D(\A_DOUT_TEMPR63[13] ), .Y(
        OR4_2175_Y));
    OR4 OR4_961 (.A(\A_DOUT_TEMPR95[38] ), .B(\A_DOUT_TEMPR96[38] ), 
        .C(\A_DOUT_TEMPR97[38] ), .D(\A_DOUT_TEMPR98[38] ), .Y(
        OR4_961_Y));
    OR2 OR2_71 (.A(\A_DOUT_TEMPR72[29] ), .B(\A_DOUT_TEMPR73[29] ), .Y(
        OR2_71_Y));
    OR4 OR4_1422 (.A(OR4_353_Y), .B(OR4_1251_Y), .C(OR4_415_Y), .D(
        OR4_2375_Y), .Y(OR4_1422_Y));
    OR4 OR4_1053 (.A(OR4_251_Y), .B(OR4_1812_Y), .C(OR4_2660_Y), .D(
        OR4_1664_Y), .Y(OR4_1053_Y));
    CFG2 #( .INIT(4'h8) )  \AND2WBYTEENA[4]  (.A(A_WBYTE_EN[2]), .B(
        A_WEN), .Y(\WBYTEENA[4] ));
    OR4 OR4_2019 (.A(\B_DOUT_TEMPR75[22] ), .B(\B_DOUT_TEMPR76[22] ), 
        .C(\B_DOUT_TEMPR77[22] ), .D(\B_DOUT_TEMPR78[22] ), .Y(
        OR4_2019_Y));
    OR4 OR4_2854 (.A(\B_DOUT_TEMPR16[29] ), .B(\B_DOUT_TEMPR17[29] ), 
        .C(\B_DOUT_TEMPR18[29] ), .D(\B_DOUT_TEMPR19[29] ), .Y(
        OR4_2854_Y));
    OR4 OR4_2704 (.A(\B_DOUT_TEMPR4[24] ), .B(\B_DOUT_TEMPR5[24] ), .C(
        \B_DOUT_TEMPR6[24] ), .D(\B_DOUT_TEMPR7[24] ), .Y(OR4_2704_Y));
    OR4 OR4_1103 (.A(OR4_2513_Y), .B(OR4_2224_Y), .C(OR4_2261_Y), .D(
        OR4_1856_Y), .Y(OR4_1103_Y));
    OR4 OR4_1428 (.A(\B_DOUT_TEMPR99[14] ), .B(\B_DOUT_TEMPR100[14] ), 
        .C(\B_DOUT_TEMPR101[14] ), .D(\B_DOUT_TEMPR102[14] ), .Y(
        OR4_1428_Y));
    OR4 OR4_1651 (.A(\B_DOUT_TEMPR115[21] ), .B(\B_DOUT_TEMPR116[21] ), 
        .C(\B_DOUT_TEMPR117[21] ), .D(\B_DOUT_TEMPR118[21] ), .Y(
        OR4_1651_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%112%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R112C4 (
        .A_DOUT({nc28140, nc28141, nc28142, nc28143, nc28144, nc28145, 
        nc28146, nc28147, nc28148, nc28149, nc28150, nc28151, nc28152, 
        nc28153, nc28154, \A_DOUT_TEMPR112[24] , \A_DOUT_TEMPR112[23] , 
        \A_DOUT_TEMPR112[22] , \A_DOUT_TEMPR112[21] , 
        \A_DOUT_TEMPR112[20] }), .B_DOUT({nc28155, nc28156, nc28157, 
        nc28158, nc28159, nc28160, nc28161, nc28162, nc28163, nc28164, 
        nc28165, nc28166, nc28167, nc28168, nc28169, 
        \B_DOUT_TEMPR112[24] , \B_DOUT_TEMPR112[23] , 
        \B_DOUT_TEMPR112[22] , \B_DOUT_TEMPR112[21] , 
        \B_DOUT_TEMPR112[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[112][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 \OR4_B_DOUT[15]  (.A(OR4_2084_Y), .B(OR4_2299_Y), .C(OR4_71_Y), 
        .D(OR4_899_Y), .Y(B_DOUT[15]));
    OR4 OR4_659 (.A(\A_DOUT_TEMPR60[16] ), .B(\A_DOUT_TEMPR61[16] ), 
        .C(\A_DOUT_TEMPR62[16] ), .D(\A_DOUT_TEMPR63[16] ), .Y(
        OR4_659_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%88%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R88C3 (
        .A_DOUT({nc28170, nc28171, nc28172, nc28173, nc28174, nc28175, 
        nc28176, nc28177, nc28178, nc28179, nc28180, nc28181, nc28182, 
        nc28183, nc28184, \A_DOUT_TEMPR88[19] , \A_DOUT_TEMPR88[18] , 
        \A_DOUT_TEMPR88[17] , \A_DOUT_TEMPR88[16] , 
        \A_DOUT_TEMPR88[15] }), .B_DOUT({nc28185, nc28186, nc28187, 
        nc28188, nc28189, nc28190, nc28191, nc28192, nc28193, nc28194, 
        nc28195, nc28196, nc28197, nc28198, nc28199, 
        \B_DOUT_TEMPR88[19] , \B_DOUT_TEMPR88[18] , 
        \B_DOUT_TEMPR88[17] , \B_DOUT_TEMPR88[16] , 
        \B_DOUT_TEMPR88[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[88][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2519 (.A(\A_DOUT_TEMPR111[33] ), .B(\A_DOUT_TEMPR112[33] ), 
        .C(\A_DOUT_TEMPR113[33] ), .D(\A_DOUT_TEMPR114[33] ), .Y(
        OR4_2519_Y));
    OR4 OR4_1878 (.A(OR4_13_Y), .B(OR4_2534_Y), .C(OR4_171_Y), .D(
        OR4_487_Y), .Y(OR4_1878_Y));
    OR4 OR4_2401 (.A(OR4_979_Y), .B(OR4_1764_Y), .C(OR4_840_Y), .D(
        OR4_529_Y), .Y(OR4_2401_Y));
    OR4 OR4_476 (.A(\A_DOUT_TEMPR56[14] ), .B(\A_DOUT_TEMPR57[14] ), 
        .C(\A_DOUT_TEMPR58[14] ), .D(\A_DOUT_TEMPR59[14] ), .Y(
        OR4_476_Y));
    OR4 OR4_1753 (.A(\A_DOUT_TEMPR87[39] ), .B(\A_DOUT_TEMPR88[39] ), 
        .C(\A_DOUT_TEMPR89[39] ), .D(\A_DOUT_TEMPR90[39] ), .Y(
        OR4_1753_Y));
    OR4 OR4_1002 (.A(\B_DOUT_TEMPR16[9] ), .B(\B_DOUT_TEMPR17[9] ), .C(
        \B_DOUT_TEMPR18[9] ), .D(\B_DOUT_TEMPR19[9] ), .Y(OR4_1002_Y));
    OR4 OR4_1947 (.A(\A_DOUT_TEMPR32[37] ), .B(\A_DOUT_TEMPR33[37] ), 
        .C(\A_DOUT_TEMPR34[37] ), .D(\A_DOUT_TEMPR35[37] ), .Y(
        OR4_1947_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%84%1%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R84C1 (
        .A_DOUT({nc28200, nc28201, nc28202, nc28203, nc28204, nc28205, 
        nc28206, nc28207, nc28208, nc28209, nc28210, nc28211, nc28212, 
        nc28213, nc28214, \A_DOUT_TEMPR84[9] , \A_DOUT_TEMPR84[8] , 
        \A_DOUT_TEMPR84[7] , \A_DOUT_TEMPR84[6] , \A_DOUT_TEMPR84[5] })
        , .B_DOUT({nc28215, nc28216, nc28217, nc28218, nc28219, 
        nc28220, nc28221, nc28222, nc28223, nc28224, nc28225, nc28226, 
        nc28227, nc28228, nc28229, \B_DOUT_TEMPR84[9] , 
        \B_DOUT_TEMPR84[8] , \B_DOUT_TEMPR84[7] , \B_DOUT_TEMPR84[6] , 
        \B_DOUT_TEMPR84[5] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[84][1] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[9], 
        A_DIN[8], A_DIN[7], A_DIN[6], A_DIN[5]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[2] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[21] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[9], B_DIN[8], 
        B_DIN[7], B_DIN[6], B_DIN[5]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[2] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2071 (.A(OR4_2282_Y), .B(OR4_2695_Y), .C(OR4_385_Y), .D(
        OR4_1225_Y), .Y(OR4_2071_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%80%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R80C4 (
        .A_DOUT({nc28230, nc28231, nc28232, nc28233, nc28234, nc28235, 
        nc28236, nc28237, nc28238, nc28239, nc28240, nc28241, nc28242, 
        nc28243, nc28244, \A_DOUT_TEMPR80[24] , \A_DOUT_TEMPR80[23] , 
        \A_DOUT_TEMPR80[22] , \A_DOUT_TEMPR80[21] , 
        \A_DOUT_TEMPR80[20] }), .B_DOUT({nc28245, nc28246, nc28247, 
        nc28248, nc28249, nc28250, nc28251, nc28252, nc28253, nc28254, 
        nc28255, nc28256, nc28257, nc28258, nc28259, 
        \B_DOUT_TEMPR80[24] , \B_DOUT_TEMPR80[23] , 
        \B_DOUT_TEMPR80[22] , \B_DOUT_TEMPR80[21] , 
        \B_DOUT_TEMPR80[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[80][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1155 (.A(OR4_1357_Y), .B(OR4_2389_Y), .C(OR4_847_Y), .D(
        OR4_2390_Y), .Y(OR4_1155_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%100%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R100C4 (
        .A_DOUT({nc28260, nc28261, nc28262, nc28263, nc28264, nc28265, 
        nc28266, nc28267, nc28268, nc28269, nc28270, nc28271, nc28272, 
        nc28273, nc28274, \A_DOUT_TEMPR100[24] , \A_DOUT_TEMPR100[23] , 
        \A_DOUT_TEMPR100[22] , \A_DOUT_TEMPR100[21] , 
        \A_DOUT_TEMPR100[20] }), .B_DOUT({nc28275, nc28276, nc28277, 
        nc28278, nc28279, nc28280, nc28281, nc28282, nc28283, nc28284, 
        nc28285, nc28286, nc28287, nc28288, nc28289, 
        \B_DOUT_TEMPR100[24] , \B_DOUT_TEMPR100[23] , 
        \B_DOUT_TEMPR100[22] , \B_DOUT_TEMPR100[21] , 
        \B_DOUT_TEMPR100[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[100][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , \BLKY1[0] , \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2788 (.A(\A_DOUT_TEMPR103[33] ), .B(\A_DOUT_TEMPR104[33] ), 
        .C(\A_DOUT_TEMPR105[33] ), .D(\A_DOUT_TEMPR106[33] ), .Y(
        OR4_2788_Y));
    OR4 OR4_2312 (.A(\A_DOUT_TEMPR36[13] ), .B(\A_DOUT_TEMPR37[13] ), 
        .C(\A_DOUT_TEMPR38[13] ), .D(\A_DOUT_TEMPR39[13] ), .Y(
        OR4_2312_Y));
    OR4 OR4_889 (.A(\B_DOUT_TEMPR36[35] ), .B(\B_DOUT_TEMPR37[35] ), 
        .C(\B_DOUT_TEMPR38[35] ), .D(\B_DOUT_TEMPR39[35] ), .Y(
        OR4_889_Y));
    OR4 OR4_953 (.A(\A_DOUT_TEMPR20[20] ), .B(\A_DOUT_TEMPR21[20] ), 
        .C(\A_DOUT_TEMPR22[20] ), .D(\A_DOUT_TEMPR23[20] ), .Y(
        OR4_953_Y));
    OR4 OR4_1520 (.A(\A_DOUT_TEMPR107[13] ), .B(\A_DOUT_TEMPR108[13] ), 
        .C(\A_DOUT_TEMPR109[13] ), .D(\A_DOUT_TEMPR110[13] ), .Y(
        OR4_1520_Y));
    OR4 OR4_2943 (.A(\A_DOUT_TEMPR87[32] ), .B(\A_DOUT_TEMPR88[32] ), 
        .C(\A_DOUT_TEMPR89[32] ), .D(\A_DOUT_TEMPR90[32] ), .Y(
        OR4_2943_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%102%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R102C3 (
        .A_DOUT({nc28290, nc28291, nc28292, nc28293, nc28294, nc28295, 
        nc28296, nc28297, nc28298, nc28299, nc28300, nc28301, nc28302, 
        nc28303, nc28304, \A_DOUT_TEMPR102[19] , \A_DOUT_TEMPR102[18] , 
        \A_DOUT_TEMPR102[17] , \A_DOUT_TEMPR102[16] , 
        \A_DOUT_TEMPR102[15] }), .B_DOUT({nc28305, nc28306, nc28307, 
        nc28308, nc28309, nc28310, nc28311, nc28312, nc28313, nc28314, 
        nc28315, nc28316, nc28317, nc28318, nc28319, 
        \B_DOUT_TEMPR102[19] , \B_DOUT_TEMPR102[18] , 
        \B_DOUT_TEMPR102[17] , \B_DOUT_TEMPR102[16] , 
        \B_DOUT_TEMPR102[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[102][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[25] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[25] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], 
        B_DIN[17], B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%61%5%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R61C5 (
        .A_DOUT({nc28320, nc28321, nc28322, nc28323, nc28324, nc28325, 
        nc28326, nc28327, nc28328, nc28329, nc28330, nc28331, nc28332, 
        nc28333, nc28334, \A_DOUT_TEMPR61[29] , \A_DOUT_TEMPR61[28] , 
        \A_DOUT_TEMPR61[27] , \A_DOUT_TEMPR61[26] , 
        \A_DOUT_TEMPR61[25] }), .B_DOUT({nc28335, nc28336, nc28337, 
        nc28338, nc28339, nc28340, nc28341, nc28342, nc28343, nc28344, 
        nc28345, nc28346, nc28347, nc28348, nc28349, 
        \B_DOUT_TEMPR61[29] , \B_DOUT_TEMPR61[28] , 
        \B_DOUT_TEMPR61[27] , \B_DOUT_TEMPR61[26] , 
        \B_DOUT_TEMPR61[25] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[61][5] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[29], 
        A_DIN[28], A_DIN[27], A_DIN[26], A_DIN[25]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[10] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[15] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[29], B_DIN[28], 
        B_DIN[27], B_DIN[26], B_DIN[25]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[10] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_281 (.A(OR4_2050_Y), .B(OR4_427_Y), .C(OR4_2981_Y), .D(
        OR4_2658_Y), .Y(OR4_281_Y));
    OR4 OR4_2 (.A(OR4_482_Y), .B(OR4_1393_Y), .C(OR4_2022_Y), .D(
        OR4_1228_Y), .Y(OR4_2_Y));
    OR4 OR4_881 (.A(\B_DOUT_TEMPR60[10] ), .B(\B_DOUT_TEMPR61[10] ), 
        .C(\B_DOUT_TEMPR62[10] ), .D(\B_DOUT_TEMPR63[10] ), .Y(
        OR4_881_Y));
    OR4 OR4_99 (.A(\A_DOUT_TEMPR44[27] ), .B(\A_DOUT_TEMPR45[27] ), .C(
        \A_DOUT_TEMPR46[27] ), .D(\A_DOUT_TEMPR47[27] ), .Y(OR4_99_Y));
    OR4 OR4_1460 (.A(\A_DOUT_TEMPR28[15] ), .B(\A_DOUT_TEMPR29[15] ), 
        .C(\A_DOUT_TEMPR30[15] ), .D(\A_DOUT_TEMPR31[15] ), .Y(
        OR4_1460_Y));
    OR4 OR4_1499 (.A(\B_DOUT_TEMPR12[8] ), .B(\B_DOUT_TEMPR13[8] ), .C(
        \B_DOUT_TEMPR14[8] ), .D(\B_DOUT_TEMPR15[8] ), .Y(OR4_1499_Y));
    OR4 OR4_1051 (.A(\B_DOUT_TEMPR56[7] ), .B(\B_DOUT_TEMPR57[7] ), .C(
        \B_DOUT_TEMPR58[7] ), .D(\B_DOUT_TEMPR59[7] ), .Y(OR4_1051_Y));
    OR4 OR4_964 (.A(\B_DOUT_TEMPR0[2] ), .B(\B_DOUT_TEMPR1[2] ), .C(
        \B_DOUT_TEMPR2[2] ), .D(\B_DOUT_TEMPR3[2] ), .Y(OR4_964_Y));
    OR4 OR4_1840 (.A(\B_DOUT_TEMPR111[21] ), .B(\B_DOUT_TEMPR112[21] ), 
        .C(\B_DOUT_TEMPR113[21] ), .D(\B_DOUT_TEMPR114[21] ), .Y(
        OR4_1840_Y));
    OR4 OR4_68 (.A(\B_DOUT_TEMPR40[27] ), .B(\B_DOUT_TEMPR41[27] ), .C(
        \B_DOUT_TEMPR42[27] ), .D(\B_DOUT_TEMPR43[27] ), .Y(OR4_68_Y));
    OR4 OR4_419 (.A(\B_DOUT_TEMPR12[4] ), .B(\B_DOUT_TEMPR13[4] ), .C(
        \B_DOUT_TEMPR14[4] ), .D(\B_DOUT_TEMPR15[4] ), .Y(OR4_419_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%77%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R77C4 (
        .A_DOUT({nc28350, nc28351, nc28352, nc28353, nc28354, nc28355, 
        nc28356, nc28357, nc28358, nc28359, nc28360, nc28361, nc28362, 
        nc28363, nc28364, \A_DOUT_TEMPR77[24] , \A_DOUT_TEMPR77[23] , 
        \A_DOUT_TEMPR77[22] , \A_DOUT_TEMPR77[21] , 
        \A_DOUT_TEMPR77[20] }), .B_DOUT({nc28365, nc28366, nc28367, 
        nc28368, nc28369, nc28370, nc28371, nc28372, nc28373, nc28374, 
        nc28375, nc28376, nc28377, nc28378, nc28379, 
        \B_DOUT_TEMPR77[24] , \B_DOUT_TEMPR77[23] , 
        \B_DOUT_TEMPR77[22] , \B_DOUT_TEMPR77[21] , 
        \B_DOUT_TEMPR77[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[77][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[19] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2904 (.A(\B_DOUT_TEMPR107[1] ), .B(\B_DOUT_TEMPR108[1] ), 
        .C(\B_DOUT_TEMPR109[1] ), .D(\B_DOUT_TEMPR110[1] ), .Y(
        OR4_2904_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%98%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R98C6 (
        .A_DOUT({nc28380, nc28381, nc28382, nc28383, nc28384, nc28385, 
        nc28386, nc28387, nc28388, nc28389, nc28390, nc28391, nc28392, 
        nc28393, nc28394, \A_DOUT_TEMPR98[34] , \A_DOUT_TEMPR98[33] , 
        \A_DOUT_TEMPR98[32] , \A_DOUT_TEMPR98[31] , 
        \A_DOUT_TEMPR98[30] }), .B_DOUT({nc28395, nc28396, nc28397, 
        nc28398, nc28399, nc28400, nc28401, nc28402, nc28403, nc28404, 
        nc28405, nc28406, nc28407, nc28408, nc28409, 
        \B_DOUT_TEMPR98[34] , \B_DOUT_TEMPR98[33] , 
        \B_DOUT_TEMPR98[32] , \B_DOUT_TEMPR98[31] , 
        \B_DOUT_TEMPR98[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[98][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[24] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[24] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2341 (.A(OR4_2072_Y), .B(OR4_1405_Y), .C(OR2_5_Y), .D(
        \B_DOUT_TEMPR74[7] ), .Y(OR4_2341_Y));
    OR4 OR4_75 (.A(OR4_2852_Y), .B(OR4_298_Y), .C(OR4_1789_Y), .D(
        OR4_301_Y), .Y(OR4_75_Y));
    OR4 OR4_3037 (.A(\B_DOUT_TEMPR40[5] ), .B(\B_DOUT_TEMPR41[5] ), .C(
        \B_DOUT_TEMPR42[5] ), .D(\B_DOUT_TEMPR43[5] ), .Y(OR4_3037_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%115%4%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R115C4 (
        .A_DOUT({nc28410, nc28411, nc28412, nc28413, nc28414, nc28415, 
        nc28416, nc28417, nc28418, nc28419, nc28420, nc28421, nc28422, 
        nc28423, nc28424, \A_DOUT_TEMPR115[24] , \A_DOUT_TEMPR115[23] , 
        \A_DOUT_TEMPR115[22] , \A_DOUT_TEMPR115[21] , 
        \A_DOUT_TEMPR115[20] }), .B_DOUT({nc28425, nc28426, nc28427, 
        nc28428, nc28429, nc28430, nc28431, nc28432, nc28433, nc28434, 
        nc28435, nc28436, nc28437, nc28438, nc28439, 
        \B_DOUT_TEMPR115[24] , \B_DOUT_TEMPR115[23] , 
        \B_DOUT_TEMPR115[22] , \B_DOUT_TEMPR115[21] , 
        \B_DOUT_TEMPR115[20] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[115][4] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[28] , A_ADDR[13], 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[24], 
        A_DIN[23], A_DIN[22], A_DIN[21], A_DIN[20]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[8] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[28] , B_ADDR[13], B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[24], B_DIN[23], 
        B_DIN[22], B_DIN[21], B_DIN[20]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[8] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%36%3%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R36C3 (
        .A_DOUT({nc28440, nc28441, nc28442, nc28443, nc28444, nc28445, 
        nc28446, nc28447, nc28448, nc28449, nc28450, nc28451, nc28452, 
        nc28453, nc28454, \A_DOUT_TEMPR36[19] , \A_DOUT_TEMPR36[18] , 
        \A_DOUT_TEMPR36[17] , \A_DOUT_TEMPR36[16] , 
        \A_DOUT_TEMPR36[15] }), .B_DOUT({nc28455, nc28456, nc28457, 
        nc28458, nc28459, nc28460, nc28461, nc28462, nc28463, nc28464, 
        nc28465, nc28466, nc28467, nc28468, nc28469, 
        \B_DOUT_TEMPR36[19] , \B_DOUT_TEMPR36[18] , 
        \B_DOUT_TEMPR36[17] , \B_DOUT_TEMPR36[16] , 
        \B_DOUT_TEMPR36[15] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[36][3] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[19], 
        A_DIN[18], A_DIN[17], A_DIN[16], A_DIN[15]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[6] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[19], B_DIN[18], B_DIN[17], 
        B_DIN[16], B_DIN[15]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[6] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_2906 (.A(\B_DOUT_TEMPR68[35] ), .B(\B_DOUT_TEMPR69[35] ), 
        .C(\B_DOUT_TEMPR70[35] ), .D(\B_DOUT_TEMPR71[35] ), .Y(
        OR4_2906_Y));
    OR4 OR4_2841 (.A(OR4_2003_Y), .B(OR4_527_Y), .C(OR4_1369_Y), .D(
        OR4_377_Y), .Y(OR4_2841_Y));
    OR4 OR4_1844 (.A(OR4_2446_Y), .B(OR4_1773_Y), .C(OR4_985_Y), .D(
        OR4_2960_Y), .Y(OR4_1844_Y));
    OR4 OR4_827 (.A(\B_DOUT_TEMPR95[32] ), .B(\B_DOUT_TEMPR96[32] ), 
        .C(\B_DOUT_TEMPR97[32] ), .D(\B_DOUT_TEMPR98[32] ), .Y(
        OR4_827_Y));
    OR4 OR4_406 (.A(\B_DOUT_TEMPR111[19] ), .B(\B_DOUT_TEMPR112[19] ), 
        .C(\B_DOUT_TEMPR113[19] ), .D(\B_DOUT_TEMPR114[19] ), .Y(
        OR4_406_Y));
    OR4 OR4_1265 (.A(\A_DOUT_TEMPR115[7] ), .B(\A_DOUT_TEMPR116[7] ), 
        .C(\A_DOUT_TEMPR117[7] ), .D(\A_DOUT_TEMPR118[7] ), .Y(
        OR4_1265_Y));
    OR4 OR4_1778 (.A(\B_DOUT_TEMPR95[5] ), .B(\B_DOUT_TEMPR96[5] ), .C(
        \B_DOUT_TEMPR97[5] ), .D(\B_DOUT_TEMPR98[5] ), .Y(OR4_1778_Y));
    OR4 OR4_2515 (.A(\A_DOUT_TEMPR64[3] ), .B(\A_DOUT_TEMPR65[3] ), .C(
        \A_DOUT_TEMPR66[3] ), .D(\A_DOUT_TEMPR67[3] ), .Y(OR4_2515_Y));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%26%0%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R26C0 (
        .A_DOUT({nc28470, nc28471, nc28472, nc28473, nc28474, nc28475, 
        nc28476, nc28477, nc28478, nc28479, nc28480, nc28481, nc28482, 
        nc28483, nc28484, \A_DOUT_TEMPR26[4] , \A_DOUT_TEMPR26[3] , 
        \A_DOUT_TEMPR26[2] , \A_DOUT_TEMPR26[1] , \A_DOUT_TEMPR26[0] })
        , .B_DOUT({nc28485, nc28486, nc28487, nc28488, nc28489, 
        nc28490, nc28491, nc28492, nc28493, nc28494, nc28495, nc28496, 
        nc28497, nc28498, nc28499, \B_DOUT_TEMPR26[4] , 
        \B_DOUT_TEMPR26[3] , \B_DOUT_TEMPR26[2] , \B_DOUT_TEMPR26[1] , 
        \B_DOUT_TEMPR26[0] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[26][0] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[6] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[4], 
        A_DIN[3], A_DIN[2], A_DIN[1], A_DIN[0]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[0] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[6] , B_ADDR[13], \BLKY0[0] }), .B_CLK(
        B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, B_DIN[4], B_DIN[3], B_DIN[2], 
        B_DIN[1], B_DIN[0]}), .B_REN(VCC), .B_WEN({GND, \WBYTEENB[0] })
        , .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), 
        .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({GND, VCC, GND}), 
        .A_WMODE({GND, GND}), .A_BYPASS(VCC), .B_WIDTH({GND, VCC, GND})
        , .B_WMODE({GND, GND}), .B_BYPASS(VCC), .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%42%7%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R42C7 (
        .A_DOUT({nc28500, nc28501, nc28502, nc28503, nc28504, nc28505, 
        nc28506, nc28507, nc28508, nc28509, nc28510, nc28511, nc28512, 
        nc28513, nc28514, \A_DOUT_TEMPR42[39] , \A_DOUT_TEMPR42[38] , 
        \A_DOUT_TEMPR42[37] , \A_DOUT_TEMPR42[36] , 
        \A_DOUT_TEMPR42[35] }), .B_DOUT({nc28515, nc28516, nc28517, 
        nc28518, nc28519, nc28520, nc28521, nc28522, nc28523, nc28524, 
        nc28525, nc28526, nc28527, nc28528, nc28529, 
        \B_DOUT_TEMPR42[39] , \B_DOUT_TEMPR42[38] , 
        \B_DOUT_TEMPR42[37] , \B_DOUT_TEMPR42[36] , 
        \B_DOUT_TEMPR42[35] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[42][7] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[10] , A_ADDR[13], 
        \BLKX0[0] }), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[39], 
        A_DIN[38], A_DIN[37], A_DIN[36], A_DIN[35]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[14] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[10] , B_ADDR[13], \BLKY0[0] }), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[39], B_DIN[38], 
        B_DIN[37], B_DIN[36], B_DIN[35]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[14] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    RAM1K20 #( .RAMINDEX("PF_SRAM_AHBL_AXI_C0%487424-487424%40-40%POWER%73%6%DUAL-PORT%ECC_EN-0")
         )  PF_SRAM_AHBL_AXI_C0_PF_DPSRAM_AHB_AXI_0_PF_DPSRAM_R73C6 (
        .A_DOUT({nc28530, nc28531, nc28532, nc28533, nc28534, nc28535, 
        nc28536, nc28537, nc28538, nc28539, nc28540, nc28541, nc28542, 
        nc28543, nc28544, \A_DOUT_TEMPR73[34] , \A_DOUT_TEMPR73[33] , 
        \A_DOUT_TEMPR73[32] , \A_DOUT_TEMPR73[31] , 
        \A_DOUT_TEMPR73[30] }), .B_DOUT({nc28545, nc28546, nc28547, 
        nc28548, nc28549, nc28550, nc28551, nc28552, nc28553, nc28554, 
        nc28555, nc28556, nc28557, nc28558, nc28559, 
        \B_DOUT_TEMPR73[34] , \B_DOUT_TEMPR73[33] , 
        \B_DOUT_TEMPR73[32] , \B_DOUT_TEMPR73[31] , 
        \B_DOUT_TEMPR73[30] }), .DB_DETECT(), .SB_CORRECT(), 
        .ACCESS_BUSY(\ACCESS_BUSY[73][6] ), .A_ADDR({A_ADDR[11], 
        A_ADDR[10], A_ADDR[9], A_ADDR[8], A_ADDR[7], A_ADDR[6], 
        A_ADDR[5], A_ADDR[4], A_ADDR[3], A_ADDR[2], A_ADDR[1], 
        A_ADDR[0], GND, GND}), .A_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        A_ADDR[12]}), .A_CLK(A_CLK), .A_DIN({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, A_DIN[34], 
        A_DIN[33], A_DIN[32], A_DIN[31], A_DIN[30]}), .A_REN(A_REN), 
        .A_WEN({GND, \WBYTEENA[12] }), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(
        VCC), .A_DOUT_SRST_N(VCC), .B_ADDR({B_ADDR[11], B_ADDR[10], 
        B_ADDR[9], B_ADDR[8], B_ADDR[7], B_ADDR[6], B_ADDR[5], 
        B_ADDR[4], B_ADDR[3], B_ADDR[2], B_ADDR[1], B_ADDR[0], GND, 
        GND}), .B_BLK_EN({\BLKY2[18] , \BLKY1[0] , B_ADDR[12]}), 
        .B_CLK(B_CLK), .B_DIN({GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, B_DIN[34], B_DIN[33], 
        B_DIN[32], B_DIN[31], B_DIN[30]}), .B_REN(VCC), .B_WEN({GND, 
        \WBYTEENB[12] }), .B_DOUT_EN(VCC), .B_DOUT_ARST_N(VCC), 
        .B_DOUT_SRST_N(VCC), .ECC_EN(GND), .BUSY_FB(GND), .A_WIDTH({
        GND, VCC, GND}), .A_WMODE({GND, GND}), .A_BYPASS(VCC), 
        .B_WIDTH({GND, VCC, GND}), .B_WMODE({GND, GND}), .B_BYPASS(VCC)
        , .ECC_BYPASS(GND));
    OR4 OR4_1315 (.A(OR4_416_Y), .B(OR4_2473_Y), .C(OR4_2698_Y), .D(
        OR4_2486_Y), .Y(OR4_1315_Y));
    OR4 OR4_1390 (.A(\A_DOUT_TEMPR75[16] ), .B(\A_DOUT_TEMPR76[16] ), 
        .C(\A_DOUT_TEMPR77[16] ), .D(\A_DOUT_TEMPR78[16] ), .Y(
        OR4_1390_Y));
    OR4 OR4_1497 (.A(\A_DOUT_TEMPR56[34] ), .B(\A_DOUT_TEMPR57[34] ), 
        .C(\A_DOUT_TEMPR58[34] ), .D(\A_DOUT_TEMPR59[34] ), .Y(
        OR4_1497_Y));
    OR4 OR4_1925 (.A(\B_DOUT_TEMPR20[22] ), .B(\B_DOUT_TEMPR21[22] ), 
        .C(\B_DOUT_TEMPR22[22] ), .D(\B_DOUT_TEMPR23[22] ), .Y(
        OR4_1925_Y));
    OR4 OR4_111 (.A(\B_DOUT_TEMPR87[5] ), .B(\B_DOUT_TEMPR88[5] ), .C(
        \B_DOUT_TEMPR89[5] ), .D(\B_DOUT_TEMPR90[5] ), .Y(OR4_111_Y));
    OR4 OR4_2532 (.A(\B_DOUT_TEMPR95[2] ), .B(\B_DOUT_TEMPR96[2] ), .C(
        \B_DOUT_TEMPR97[2] ), .D(\B_DOUT_TEMPR98[2] ), .Y(OR4_2532_Y));
    OR4 OR4_438 (.A(\A_DOUT_TEMPR103[31] ), .B(\A_DOUT_TEMPR104[31] ), 
        .C(\A_DOUT_TEMPR105[31] ), .D(\A_DOUT_TEMPR106[31] ), .Y(
        OR4_438_Y));
    OR4 OR4_2868 (.A(OR4_2341_Y), .B(OR4_2331_Y), .C(OR4_1524_Y), .D(
        OR4_461_Y), .Y(OR4_2868_Y));
    OR2 OR2_47 (.A(\B_DOUT_TEMPR72[4] ), .B(\B_DOUT_TEMPR73[4] ), .Y(
        OR2_47_Y));
    OR4 OR4_534 (.A(\B_DOUT_TEMPR28[2] ), .B(\B_DOUT_TEMPR29[2] ), .C(
        \B_DOUT_TEMPR30[2] ), .D(\B_DOUT_TEMPR31[2] ), .Y(OR4_534_Y));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
